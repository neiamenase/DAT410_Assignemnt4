jag förklarar europaparlamentets session återupptagen efter avbrottet den 17 december . jag vill på nytt önska er ett gott nytt år och jag hoppas att ni haft en trevlig semester .
som ni kunnat konstatera ägde &quot; den stora år 2000-buggen &quot; aldrig rum . däremot har invånarna i ett antal av våra medlemsländer drabbats av naturkatastrofer som verkligen varit förskräckliga .
ni har begärt en debatt i ämnet under sammanträdesperiodens kommande dagar .
till dess vill jag att vi , som ett antal kolleger begärt , håller en tyst minut för offren för bl.a. stormarna i de länder i europeiska unionen som drabbats .
jag ber er resa er för en tyst minut .
ni känner till från media att det skett en rad bombexplosioner och mord i sri lanka .
en av de personer som mycket nyligen mördades i sri lanka var kumar ponnambalam , som besökte europaparlamentet för bara några månader sedan .
skulle det vara möjligt för er , fru talman , att skriva ett brev till den srilankesiska presidenten i vilket parlamentets beklagande uttrycks över hans och de övriga brutala dödsfallen i sri lanka och uppmanar henne att göra allt som står i hennes makt för att få en fredlig lösning på en mycket komplicerad situation ?
ja , herr evans , jag tror att ett initiativ i den riktning ni just föreslagit skulle vara mycket lämpligt .
om kammaren instämmer skall jag göra som herr evans föreslagit .
jag skulle vilja ha råd från er vad gäller artikel 143 om avvisning av ett ärende som otillåtligt .
min fråga har att göra med något som kommer att behandlas på torsdag och som jag då kommer att ta upp igen .
cunhas betänkande om de fleråriga utvecklingsprogrammen behandlas i parlamentet på torsdag och det innehåller ett förslag i punkt 6 om att något slag av kvoteringspåföljder bör införas för länder som misslyckas med att uppfylla sina årliga mål rörande minskning av flottorna .
i betänkandet står det att detta bör göras trots principen om relativ stabilitet .
jag anser att principen om relativ stabilitet är en grundläggande rättsprincip inom den gemensamma fiskeripolitiken , och ett förslag som skulle undergräva den måste betraktas som rättsligt otillåtligt .
jag vill veta om jag kan göra en sådan invändning mot ett betänkande , som alltså inte är ett lagförslag , och om det är något som jag har behörighet att göra på torsdag .
det är faktiskt just vid det tillfället som ni , om ni vill , kan ta upp denna fråga , dvs. på torsdag innan betänkandet läggs fram .
under årets första sammanträdesperiod för europaparlamentet bestämde man dessvärre i texas i usa att nästa torsdag avrätta en dödsdömd , en ung man på 34 år som vi kan kalla hicks .
på uppmaning av en fransk parlamentsledamot , zimeray , har redan en framställning gjorts , undertecknad av många , bland annat jag själv , men jag uppmanar er , i enlighet med de riktlinjer som europaparlamentet och hela den europeiska gemenskapen alltid har hållit fast vid , att med all den tyngd ni har i kraft av ert ämbete och den institution ni företräder , uppmana texas guvernör , bush , att uppskjuta verkställigheten och att benåda den dömde .
detta är helt i linje med de principer som vi alltid har hävdat .
tack , herr segni , det skall jag gärna göra .
det ligger faktiskt helt i linje med de ståndpunkter vårt parlament alltid antagit .
fru talman ! jag vill fästa er uppmärksamhet vid ett fall som parlamentet vid upprepade tillfällen har befattat sig med .
det gäller fallet alexander nikitin .
alla gläder vi oss åt att domstolen har friat honom och tydligt visat att tillgängligheten till miljöinformation är en konstitutionell rättighet även i ryssland .
nu är det emellertid så att han skall åtalas på nytt i och med att allmänne åklagaren överklagar .
vi är medvetna om , vilket vi också - inte minst under förra årets sista plenarsammanträde - har kunnat konstatera i en lång rad beslut , att detta inte enbart är ett juridiskt fall och att det är fel att beskylla alexander nikitin för kriminalitet och förräderi , eftersom vi som berörda parter drar nytta av de resultat han har kommit fram till .
resultaten utgör grunden för de europeiska programmen för skydd av barents hav , och därför ber jag er granska ett utkast till ett brev som skildrar de viktigaste fakta samt att i enlighet med parlamentsbesluten visa ryssland denna ståndpunkt klart och tydligt .
ja , fru schroedter , jag skall mycket gärna granska fakta rörande denna fråga när jag fått ert brev .
fru talman ! först skulle jag vilja ge er en komplimang för det faktum att ni hållit ert ord och att det nu , under det nya årets första sammanträdesperiod , faktiskt har skett en kraftig utökning av antalet tv-kanaler på våra rum .
men , fru talman , det som jag bad om har inte inträffat .
det finns nu visserligen två finska kanaler och en portugisisk , men det finns fortfarande ingen nederländsk kanal . jag bad er om en nederländsk kanal , eftersom nederländare också gärna vill ta del av nyheterna varje månad då vi blir förvisade till den här platsen .
jag skulle således på nytt vilja be er att ombesörja att vi också får en nederländsk kanal .
fru plooij-van gorsel ! jag kan tala om för er att frågan finns på föredragningslistan för kvestorernas möte på onsdag .
jag hoppas att den kommer att granskas i en positiv anda .
fru lynne ! ni har helt rätt och jag skall kontrollera om allt detta faktiskt inte har gjorts .
jag skall också överlämna problemet till kvestorerna och jag är övertygad om att de är måna om att se till att vi respekterar de regler som vi faktiskt röstat fram .
fru talman ! díez gonzález och jag har ställt några frågor angående vissa av vice ordförande de palacios åsikter som återgavs i en spansk dagstidning .
de ansvariga har inte tagit med dessa frågor på föredragningslistan , eftersom man ansåg att dessa hade besvarats vid ett tidigare sammanträde .
jag ber att man omprövar det beslutet , eftersom så inte är fallet .
de frågor som tidigare besvarats handlade om de palacios inblandning i ett särskilt ärende , inte om de uttalanden som återgavs i dagstidningen abc den 18 november i fjol .
kära kollega ! vi skall kontrollera allt detta .
jag erkänner att för närvarande förefaller saker och ting litet oklara .
vi skall alltså se över detta mycket noga så allt blir i sin ordning .
i vilket fall som helst är frågan för närvarande inte föremål för någon begäran om brådskande förfarande på torsdag .
nästa punkt på föredragningslistan är fastställande av arbetsplanen . det slutgiltiga förslaget till föredragningslista som utarbetats av talmanskonferensen vid sammanträdet den 13 januari i enlighet med artikel 110 i arbetsordningen har delats ut .
för måndag och tisdag har inga ändringar föreslagits .
beträffande onsdag :
den socialistiska gruppen har begärt att ett uttalande från kommissionen om dess strategiska mål för de fem kommande åren samt om kommissionens administrativa reform skall tas upp .
jag skulle vilja att barón crespo , som lämnat begäran , uttalar sig för att motivera den , om han vill , naturligtvis .
sedan gör vi som vi brukar : vi lyssnar till en talare för och en talare emot .
fru talman ! framläggandet av kommission prodis politiska program för hela mandatperioden bottnar i ett förslag från europeiska socialdemokratiska partiets grupp som antogs med enhällighet på talmanskonferensen i september samt ett tydligt godkännande från ordförande prodi som upprepade detta åtagande i sitt anförande i samband med tillträdandet av sitt ämbete .
detta åtagande är viktigt , med tanke på att kommissionen är det organ som enligt fördragen har ensam initiativrätt , och det utgör därför grunden till parlamentets politiska och lagstiftande verksamhet de kommande fem åren .
jag vill dessutom , fru talman , påminna om att parlamentet vid två tillfällen under föregående mandatperiod röstade om förtroendet för ordförande prodi ; man röstade på nytt om detta under denna mandatperiod i juli , och sedan , när den nya kommissionen hade påbörjat sitt arbete , gav man i september en förtroenderöst till hela kommissionen .
därför har det funnits tillräckligt mycket tid för kommissionen att förbereda sitt program och för att oss att ta del av detta och redogöra för detta inför medborgarna .
jag vill också påminna om resolutionen av den 15 september , där man rekommenderade att förslaget skulle läggas fram så snart som möjligt .
det som hände förra veckan - något som inleddes utanför talmanskonferensen , en konferens som endast utnyttjades för att bestyrka och bekräfta det beslut som fattats utanför ramarna för denna - utgör ett dilemma : antingen är det så att kommissionen inte är i stånd att presentera programmet ( i sådant fall bör den klargöra detta .
enligt ordförandens uttalanden kan man presentera programmet .
med tanke på att kommissionen företräds av vice ordförande de palacio , anser jag att vi innan omröstningen sker bör få veta huruvida kommissionen är beredd att lägga fram programmet , så som man kommit överens om ) ; annars är parlamentet inte i stånd att granska programmet , så som vissa tycks anse .
enligt min uppfattning skulle den sistnämnda hypotesen innebära att vi försummade vårt ansvar som parlament , förutom att man då skulle införa en grundtes , en okänd metod som innebär att de politiska grupperna skriftligen får ta del av kommissionens tankar kring programmet en vecka i förväg i stället för en dag i förväg , som man kommit överens om . då bör man tänka på att lagstiftningsprogrammet skall debatteras i februari , och därför skulle vi lika gärna kunna avstå från den debatten , för pressen och internet skulle redan dagen därpå tillkännage programmet för alla medborgare , och det skulle inte längre finnas någon anledning för parlamentet att ägna sig åt frågan .
eftersom min grupp anser att parlamentet är till för att lyssna , för att debattera och för att reflektera , anser vi att det inte finns något som rättfärdigar en senareläggning av debatten , och om kommissionen är beredd till det , menar vi att det fortfarande är möjligt att återupprätta det ursprungliga avtalet mellan parlamentet och kommissionen och agera på ett ansvarsfullt sätt gentemot våra medborgare .
därför innebär förslaget från europeiska socialdemokratiska partiets grupp , som fru talmannen nämnde , att kommission prodis lagstiftningsprogram läggs fram på onsdag som planerat , och att man inbegriper förslaget om en administrativ reform , för i annat fall kan en paradoxal situation uppstå : å ena sidan vägras kommissionens ordförande , med ursäkten att det inte finns något dokument , rätten att tala i parlamentet , å andra sidan omöjliggörs en debatt om reformen , eftersom parlamentet inte tidigare har fått ta del av dokumenten i fråga .
därför ber jag , fru talman , att ni uppmanar kommissionen att uttala sig och att vi därefter går till omröstning .
( applåder från pse )
jag föreslår att vi röstar om begäran från den socialistiska gruppen att på nytt föra upp kommissionens uttalande om dess strategiska mål på föredragningslistan .
beträffande onsdagen har jag också mottagit ett annat förslag beträffande den muntliga frågan om kapitalskatt .
ppe-de-gruppen begär att denna punkt skall strykas från föredragningslistan .
vill någon kollega begära ordet för gruppens räkning och motivera denna begäran ?
eftersom jag hör att det skrattas bland socialisterna : man har sagt mig att även vida kretsar inom den socialistiska gruppen gärna vill se den här punkten avförd från föredragningslistan , eftersom det vid omröstningen på talmanskonferensen saknades votum för berörda kolleger i den socialistiska arbetsgruppen .
jag vet inte huruvida denna information stämmer , men vi i ppe-de-gruppen vore i alla fall tacksamma ifall punkten ströks , då ju parlamentet redan har befattat sig med frågan flera gånger .
det finns också beslut fattade mot en sådan skatt .
därför yrkar min grupp på att punkten avförs från föredragningslistan .
tack , herr poettering .
vi skall nu lyssna till wurtz som skall uttala sig emot denna begäran .
fru talman ! jag skulle till att börja med vilja understryka poetterings bristande logik .
han har just läxat upp den socialistiska gruppen för att den ändrat sig när det gäller ett beslut som fattats med mycket liten marginal i talmanskonferensen . men han gör samma sak själv .
vi diskuterade och var eniga , utom ppe-gruppen och den liberala gruppen , och jag noterade t.o.m. , det minns ni säkert kära ordförandekolleger , att frågan inte handlar om huruvida ni är för eller emot todinskatten , utan om ni vågar höra vad kommissionen och rådet tycker om den .
jag upprepar därför förslaget att behålla denna muntliga fråga till kommissionen och rådet för att en gång för alla få veta vilken inställning dessa två instanser har till denna relativt blygsamma begäran , som ändå skulle utgöra en viktig signal till allmänheten , särskilt med tanke på den oro som uppstod efter den misslyckade konferensen i seattle .
vi skall rösta om begäran från ppe-de-gruppen som syftar till att stryka den muntliga frågan om kapitalskatt från föredragningslistan .
( parlamentet avslog begäran med 164 röster för , 166 emot . 7 ledamöter avstod från att rösta . )
fru talman ! jag skulle vilja tacka poettering för att han just gjort reklam för denna debatt .
jag undrar om även min röst har räknats , trots att den inte kunde avges på elektronisk väg , eftersom jag inte har något kort ?
jag röstade &quot; för &quot; .
om man lägger till de två kolleger som yttrat sig blir resultatet ...
fru talman ! under den tidigare omröstningen - och jag kommer att följa ert utslag i denna fråga - rörande frågan om kommissionens strategiska plan , sade jag att jag ville uttala mig före omröstningen på min grupps vägnar .
så blev inte fallet .
jag skulle uppskatta om jag vid denna punkts avslutande kunde få avge en röstförklaring på min grupps vägnar .
det skulle vara användbart för kammarens räkning att upplysa om hur folk uppfattar vad vi just gjort mot bakgrund av deras egen politiska analys .
fru talman ! jag skall inte ta upp debatten på nytt , men även jag hade begärt ordet för att ta ställning till herr barón crespos begäran .
ni lät mig aldrig komma till tals .
det beklagar jag , men omröstningen har genomförts , beslutet har fattats , alltså får det vara .
jag är ledsen , herr hänsch och herr cox , jag såg inte att ni hade begärt ordet .
jag tror ändå att ståndpunkterna är tydliga och de kommer att bekräftas i protokollet .
när vi i morgon justerar protokollet från dagens sammanträde kan de kolleger , som då anser att ståndpunkterna inte förklarats tillräckligt tydligt , begära ändringar .
jag tror att det är ett bra sätt .
naturligtvis kommer man i protokollet från morgondagens sammanträde att ta hänsyn till alla kompletterande förklaringar .
jag tror att det är bättre än att nu genomföra röstförklaringar som kommer att leda mycket långt .
vad säger ni om det , herr cox och herr hänsch ?
fru talman ! om omröstningsregistreringen på ett korrekt sätt visar hur min grupp röstade , skall jag och kan jag inte protestera mot denna .
om ert utslag innebär att jag inte kan avge en röstförklaring , accepterar jag detta men med reservation .
vi skall alltså vara mycket noggranna vid upprättandet av protokollet . det är vi för övrigt alltid .
om det inte återger ståndpunkterna tillfredsställande , kan vi eventuellt ändra i det .
( arbetsplanen fastställdes med dessa ändringar . )
säkerhetsrådgivare för transport av farligt gods
nästa punkt på föredragningslistan är andrahandsbehandlingsrekommendation ( a5-0105 / 1999 ) av koch , för utskottet för regionalpolitik , transport och turism om rådets gemensamma ståndpunkt inför europaparlamentets och rådets direktiv om harmoniseringen av examineringskraven för säkerhetsrådgivare för transport av farligt gods på väg , järnväg eller inre vattenvägar ( c5-0208 / 1999 - 1998 / 0106 ( cod ) ) .
( de ) ärade fru kommissionär , ärade fru talman , kära kolleger ! jag välkomnar utan förbehåll rådets gemensamma ståndpunkt i strävan mot att skapa en enhetlig utbildning av säkerhetsrådgivare för transport av farligt gods på landsväg , järnväg eller inre vattenvägar .
för det första : vi var tvungna att formellt börja arbeta för att kraven enligt direktiv 96 / 35 / eg skulle uppfyllas , enligt vilka medlemsländerna förpliktigas att vid hantering av farligt gods ta hjälp av ombud resp. säkerhetsrådgivare liksom att organisera utbildning , kurser och examination för dessa personer , utan att utföra detta explicit .
för det andra : genom direktivet uppnår vi a ) bättre säkerhet , såväl under transport som under omlastning av farligt gods ; b ) minskad snedvridning av konkurrensen till följd av de mest skilda nationella utbildningsstrukturer och utbildningskostnader liksom c ) lika villkor för säkerhetsrådgivare på den europeiska arbetsmarknaden .
för det tredje garanterar vi med direktivet såsom det nu föreligger som gemensam ståndpunkt , särskilt i och med att det uteslutande inskränks till miniminormer , en hög grad av flexibilitet och ringa reglering från europeiska unionens sida , och vi bidrar till stort egenansvar för medlemsländerna .
allt detta kan vi varmt välkomna i enlighet med subsidiaritetsprincipen .
jag anser att våra ändringsförslag från första behandlingen har fått vederbörlig uppmärksamhet .
de antogs , andemeningen förverkligades eller också föll de bort på grund av att aktuella europeiska bestämmelser inte infördes , t.ex. ett sanktionssystem mot överträdelser eller en komplicerad blockbildning av frågekomplex .
jag ber om samtycke till det ena enhälligt godkända ändringsförslaget från utskottet för regionalpolitik och transport , vilket gäller det tidsmässiga införlivandet av direktivet .
i och med att vi inte ger medlemsstaterna något specifikt datum för införlivandet av direktivet utan godkänner en tidsfrist på tre månader från direktivets ikraftträdande , inför vi en flexibilitetsklausul som garanterar ett omedelbart införlivande .
jag ber om samtycke .
fru talman ! vi varken kan eller får finna oss i att allt oftare höra talas om olyckor där stora skador uppstår på våra vägar , men också på järnväg eller inre vattenvägar , inte bara , men också därför att berörda personer inte tar transporten av farligt gods på tillräckligt stort allvar eller därför att okunskap eller bristande utbildning av förarna eller andra ansvariga för de olika kommunikationsmedlen alltför ofta har förvandlat en liten olycka till en stor katastrof .
jag som österrikare , men jag tror att det gäller oss alla , har fortfarande den katastrof i färskt minne som förra året kostade många människor livet i tauerntunneln , där det tog många månader av ett enormt ekonomiskt pådrag att bygga upp vad som förstördes vid branden .
den månadslånga renoveringen skar av denna viktiga trafikled mellan europas norra och södra delar .
den omväg för trafiken som detta medförde innebar för många tusen eu-medborgare en påfrestning på gränsen till det uthärdliga .
på sina håll i mitt land var det ett rent helsike .
förebyggande åtgärder måste bli vårt svar på dylika katastrofer , och med föreliggande direktivförslag skapar vi en viktig grund för att välutbildade säkerhetsrådgivare skall kunna stå till förfogande för att i tid göra det rätta .
vi får faktiskt inte nöja oss med att skapa en europeisk lag i akt och mening att skapa höjd säkerhet .
vi måste även konsekvent ge akt på att medlemsstaterna genomför våra riktlinjer inom föreskriven tidsram , och ännu viktigare , vi måste ge akt på att de sedan verkligen tillämpas också .
inte ännu ett område där vi i efterhand måste beklaga den bristande verkställigheten , tack .
jag skulle vilja ta upp en sista punkt : vi får ingalunda nöja oss med att lappa ihop ännu ett hål i säkerhetsnätet och blunda för att det återstår mycket mer att göra på området transportsäkerhet i europa .
vidare kräver jag och ber närvarande ansvarig kommissionär att så snart som möjligt lägga fram ett dokument som sörjer för bättre säkerhet i framtida tunneltrafik så att vi slipper uppleva fler katastrofer av denna vidd här i europa !
fru talman ! låt mig först och främst tacka koch för hans betänkande , i vilket han på ett mycket seriöst sätt behandlat frågan om transportsäkerhet .
han behandlar frågan om harmonisering av examineringskraven för säkerhetsrådgivare för transport av farligt gods på väg , järnväg och inre vattenvägar .
jag gratulerar honom till hans utmärkta betänkande .
transportsäkerheten har tråkigt nog diskuterats i nyheterna nyligen : tågkraschen vid paddington i london , den fruktansvärda tågkraschen i norge , de två flygkrascherna där eu-medborgare fanns ombord och naturkatastrofen utanför bretagnes kust efter erikas haveri - som alla skett inom de senaste fyra månaderna - påminner oss om att transportsäkerheten aldrig kan tas för given och de som ansvarar för att skydda allmänheten måste vara mycket motiverade och mycket kvalificerade .
föredraganden har påpekat för kammaren att rådet i sin gemensamma ståndpunkt har godkänt sex av parlamentets tio ändringsförslag som lades fram vid första behandlingen , och att andemeningen i parlamentets övriga ändringsförslag har behållits .
min grupp vill därför stödja den gemensamma ståndpunkten och ser fram emot antagandet av lagstiftningen , vilken kommer att ge oss ytterligare ett instrument i vår kamp för att göra transporterna i europeiska unionen så säkra som möjligt .
när det gäller säkerhet kommer min grupp alltid att stödja initiativ som avser att förbättra transportsäkerheten .
som händelserna under den senaste tiden visat , har vi fortfarande mycket arbete kvar på detta område .
fru talman ! i detta parlament uppmärksammas regelbundet , med rätta , hur viktig transportsäkerheten är .
de alltjämt ökande mängder gods som transporteras genom europa medför medvetet och omedvetet allehanda risker för personalen och samhällsomgivningen .
de som måste hantera dessa risker måste därför uppfylla höga krav .
de normer för detta som fastlagts i ett annat direktiv , 95 / 35 / eg , förefaller vara tillräckligt adekvata för att på ett ansvarigt sätt ge råd om hur transporter av farligt gods skall organiseras .
det gläder mig att vi också nått samförstånd med rådet i fråga om minimikraven för deras examen , även om jag hellre hade sett att enhetliga fasta normer kommit till stånd , så att examensbevisen är lika internationellt sett .
men det har visat sig att detta inte går att uppnå .
slutligen , ändringsförslaget som föredraganden föreslår är inte mer än logiskt , och därför kan jag också helhjärtat stödja detta .
herr talman , fru kommissionär , ärade kolleger ! först vill jag gratulera min kollega koch till hans betänkanden , som måhända är tekniska rapporter , men som har mycket stor betydelse för säkerheten .
jag vill endast göra några små anmärkningar .
först vill jag be fru kommissionären - och jag är övertygad om att min önskan faller i god jord - att ägna säkerhetsfrågan större uppmärksamhet , vare sig det gäller på vägar , på inre vattenvägar eller på havet .
när jag inser att den första begäran gjordes till kommissionen den 19 mars 1998 och att vi behandlar frågan här i dag - trots att parlamentet reagerade relativt snart - då tycker jag att tidsrymden är något för lång .
nu är detta inte enbart kommissionens fel , men jag tycker att vi måste reagera snabbare för att få till stånd en standardisering även här .
den andra punkten nämndes just : minimireglerna .
jag är principiellt av den åsikten att vi på många transportområden borde eftersträva ökad flexibilitet samt regelverk som gäller land för land .
när det gäller säkerheten är jag dock något skeptisk , eftersom säkerheten i låt oss säga sverige i princip inte skiljer sig från säkerheten i tyskland , italien eller österrike .
jag kan leva med dessa minimiregler , men jag ber kommissionen att verkligen uppmärksamt följa händelseutvecklingen .
om den här typen av flexibilitet i vissa länder skulle leda till bristfälliga bestämmelser , då bör vi genomföra ytterligare standardiseringar .
den tredje punkten har även den nämnts .
jag kommer ju , precis som min kollega rack , från ett transitland , där denna fråga spelar en särskild roll .
vi skall inte försämra konkurrensvillkoren ensidigt för vissa länder och förbättra dem för länder som österrike eller andra transitländer .
men jag anser att vi bör göra allt för att hålla transporten av farligt gods på så låg nivå som möjligt , och det i alla länder , transitland eller inte .
herr talman ! jag vill börja med att gratulera föredragande koch till hans utmärkta arbete och hans konstruktiva samarbete med kommissionen när det gällt att förbättra texten , föredra detta betänkande och förslag ; slutligen finns det endast ett ändringsförslag beträffande examineringskraven för säkerhetsrådgivare för transport av farligt gods på väg , järnväg eller inre vattenvägar .
vi anser att samarbetet är av stor betydelse , de gemensamma insatserna från de båda institutionerna - parlamentet och kommissionen - och samarbetet med utskottet för regionalpolitik , transport och turism , med transportgruppen närmare bestämt , fungerar alldeles utmärkt .
den gemensamma ståndpunkten inbegriper praktiskt taget alla ändringsförslag som har godkänts av kommissionen , examineringskraven för säkerhetsrådgivare har harmoniserats och , i andra behandlingen , kan vi godkänna ändringsförslaget med ett datum som är mer realistiskt än det datum som kommissionen föreslog i början , med tanke på att vi redan har debatterat den här frågan i många år .
jag vill också kort tacka de olika parlamentsledamöterna för deras insats och tala om för er , mina damer och herrar , att kommissionen prioriterar säkerheten på transportområdet .
och simpson har alldeles rätt i det han sade , att man aldrig får betrakta processen som slutförd , som avklarad eller som färdig .
processen med ett utökande av marginalerna , av säkerhetsgarantierna vid transport är en process som måste förbättras dag för dag .
i den bemärkelsen vill jag också kort ta upp problematiken med tunnlarna , som rack och swoboda hänvisade till , och som utan tvekan är en mycket känslig fråga för österrikes del , och vi måste därför bemöda oss om att förbättra säkerheten .
vid en av de större olyckor som inträffat på senare tid , var inte det transporterade godset farligt i sig .
margarin och några kilo målarfärg , som i princip inte utgjorde någon risk , kom att orsaka en riktig katastrof .
därför måste man fundera över hur man ytterligare kan skärpa de krav som garanterar en maximal säkerhet .
avslutningsvis vill jag säga att säkerheten måste iakttas vid alla typer av transporter .
den här veckan skall vi hålla en debatt där vi talar om säkerheten vid sjötransporter , till följd av katastrofen med erika , och vi kommer under det här året att få diskutera målsättningen i fråga om säkerhet vid flygtransporter .
mina damer och herrar , jag vill påpeka att säkerheten är ett mål som prioriteras av kommissionen .
och som jag kommer att säga i debatten om erika , får vi inte vänta tills det inträffar en katastrof innan vi tar itu med säkerhetsaspekten . låt oss i stället ta oss an frågan utanför sådana situationer som inte utgör annat än ett bevis på hur brådskande det är med en effektiv lösning på denna typ av problem .
jag vill än en gång rikta ett tack till alla som har medverkat och då i synnerhet föredragande koch .
transport av farligt gods på väg
nästa punkt på föredragningslistan är betänkande ( a5-0104 / 1999 ) av koch för utskottet för regionalpolitik , transport och turism om europaparlamentets och rådets direktiv om ändring av direktiv 94 / 55 / eg om tillnärmning av medlemsstaternas lagstiftning om transport av farligt gods på väg &#91; kom ( 1999 ) 158 - c5-0004 / 1999 - 1999 / 0083 ( cod ) &#93; .
) herr talman , ärade fru kommissionär , kära kolleger ! det direktiv som trädde i kraft den 1 januari 1997 om tillnärmning av medlemsstaternas lagstiftning om transport av farligt gods på väg innehåller en del övergångsbestämmelser , vars giltighet är temporär och knuten till att cen , alltså europeiska standardiseringskommittén , utarbetar bestämda regler .
de dröjsmål som har uppstått i cen : s arbete leder nu till problem med införlivandet av direktivet .
framför allt kan bilagorna inte anpassas i takt med den tekniska och industriella utvecklingen .
jag beklagar detta , för nu måste vi göra det arbete andra inte har gjort .
i så måtto accepterar jag föreliggande förslag om ändring av direktiv 94 / 55 / eg , vilket skall diskuteras i dag .
om europeiska unionen avstår från att gripa in skulle detta tvinga medlemsstaterna att ändra sina inhemska rättsliga bestämmelser för en kort period , nämligen tills cen : s arbete har slutförts , vilket drar med sig onödiga kostnader och förvirring .
den ändring av direktivet som i dag står på föredragningslistan innebär alltså ingen förändring i den standardisering av transport av farligt gods som gemenskapen har i dag .
genom denna utvidgas däremot övergångsbestämmelserna genom att gällande datum skjuts upp , de bestämmelser som inte längre är relevanta stryks och den innebär att förfarandet regleras vid a ) ad hoc-transporter av farligt gods liksom b ) införandet av mindre stränga nationella bestämmelser , särskilt vad gäller transport av mycket ringa mängder farligt gods på geografiskt sett mycket strängt avgränsade områden .
därmed ligger ändringen av direktivet helt i linje med subsidiaritetsprincipen : medlemsländerna får större befogenheter .
eu-kommissionen avgör huruvida medlemsländerna kan införa egna särskilda bestämmelser .
kommissionen stöds efter regleringsförfarandet av ett expertutskott för transport av farligt gods .
detaljerna för hur dessa befogenheter som anförtrotts kommissionen skall utövas har ändrats i rådets beslut från juni 1999 .
det förslag till ändring av direktivet gällande transport av farligt gods på väg , som skall diskuteras i dag , är dock från maj 1999 och har därför ännu inte kunnat ta hänsyn till det aktuella kommittéförfarandet .
de framlagda och av utskottet enhälligt godkända ändringsförslagen åberopar i två fall just detta förändrade kommittéförfarandet .
vi skulle vilja säkerställa att det redan i motiveringen hänvisas till detta och att den icke entydigt formulerade tidsfristen , inom vilken rådet måste fatta beslut , fastställts till högst tre månader .
därutöver hänvisas det till nödvändigheten av ökad öppenhet .
ett annat ändringsförslag tillåter medlemsländerna att införa skärpta krav , framför allt för vakuumtankar , för arbete resp. transport vid temperaturer på under minus 20 º c. detta är särskilt intressant för de nordeuropeiska regionerna .
ett sista ändringsförslag skall göra det tillåtet att fortsätta använda de tankar och tankfordon som tagits i bruk mellan den 1 januari 1997 och ikraftträdandet av detta direktiv , under förutsättning att de konstruerats och servats på vederbörligt sätt .
även om jag är medveten om att detta endast är ett litet steg mot ökad transportsäkerhet ber jag er anta betänkandet .
herr talman , bästa kolleger ! gott nytt år och gott nytt millennium !
det är första gången jag talar vid plenarsammanträdet och detta är spännande , i viss mån likt den första kärleken , men den första kärleken varade dock längre än två minuter .
jag skulle kort vilja kommentera kommissionens förslag till ändring av direktivet om transport av farligt gods på väg .
det är bra att detta direktiv utfärdas nu eftersom medlemsstaterna i annat fall skulle tvingas att ändra sina nationella bestämmelser för en mycket kort tid , en övergångsperiod , vilket i sin tur bara skulle förorsaka onödiga kostnader och än en gång öka allmänhetens grämelse över eu : s byråkrati .
i kommissionens förslag har man emellertid inte tagit hänsyn till alla aspekter , som till exempel de nordliga regionernas kalla klimat .
därför har jag föreslagit några ändringar , som godkänts i vårt utskott , till kollegan kochs i och för sig utmärkta betänkande .
mina ändringsförslag gäller köldbeständigheten hos de tankar som används för transport av dessa farliga ämnen .
enligt kommissionens förslag skulle det räcka med minus tjugo grader ; vid medelhavet har man svårt att föreställa sig att temperaturen i lappland skulle kunna sjunka betydligt lägre .
även i lappland stödjer man eu , låt oss därför även komma ihåg dem som bor där .
således föreslår jag att köldgränsen skall sänkas till minus fyrtio grader .
detta är också nödvändigt för att bibehålla nuvarande säkerhetsnivå i de nordliga områdena .
jag hoppas att mina förslag beaktas vid omröstningen i morgon .
herr talman ! tillåter ni att jag först av allt uttrycker min respekt för ert sätt att klara det flygande bytet på ordförandebänken under debatten för en stund sedan .
det var lysande .
till saken : jag anser att europas medborgare måste kunna lita på att det som transporteras på europas vägar , järnvägsnät osv. , även om det är farligt gods , transporteras så säkert som möjligt .
direktivet är ett bidrag till detta .
vad vi gör här i dag är i grund och botten ett irritationsmoment .
föredraganden koch , som vi tackar för det arbete han har utfört , har påpekat att i princip allt redan hade kunnat komma längre om det inte hade varit för försummelsen från cen , som är mycket senfärdig med att upprätta och anpassa riktlinjen .
därför kan vi bara hoppas - och denna vecka helst besluta om - att vi år 2001 äntligen får en gemensam reglering av transporten av farligt gods på väg , så att vi får en gnutta rättssäkerhet här inne och en gnutta ökad säkerhet där ute på våra vägar .
herr talman ! det betänkande som vi här behandlar innebär i sig inga stora förändringar .
de flesta av ändringsförslagen är av enbart teknisk natur .
det är dock värt att understryka att varje gång som vi fattar denna typ av beslut är det bra ur ett brett miljöperspektiv , och det är bra därför att det skapar bättre förutsättningar för den inre marknadens möjligheter att fungera .
det transporteras runtom i eu mycket stora mängder farligt gods både på vägar , järnvägar och på haven .
det gör att det är nödvändigt med ordentliga regler för hur detta skall fungera .
på område efter område får vi nu gemensamma minimiregler för medlemsländerna .
det är utomordentligt positivt , och det finns anledning att tacka föredraganden , koch , för det arbete som han har lagt ned på detta ärende .
detta är också viktigt när det gäller förutsättningarna för den inre marknaden .
om vi skall få en gemensam transportmarknad att verkligen fungera , är det viktigt , inte bara att vi har regler , utan också att dessa regler så långt som möjligt är gemensamma .
jag vill avslutningsvis gärna kommentera en tredje sak som också är väsentlig , nämligen ett ändringsförslag framlagt av ledamoten ari vatanen .
på många sätt skiljer sig förutsättningarna från ett medlemsland till ett annat .
genom att godkänna detta ändringsförslag , tar vi hänsyn till att det i de norra delarna av unionen kan vara mycket kallt .
det gör att det är nödvändigt att också ta hänsyn till hur material och förpackningar påverkas av en sådan kyla .
herr talman , det är positivt att vi i denna reglering också kan vara flexibla .
det är min förhoppning att kommissionen kan acceptera denna ändring .
herr talman ! jag vill tacka inte bara kollegan koch , utan också vice ordföranden i kommissionen för hennes klara och entydiga ställningstagande för säkerheten på transportområdet och prioriteringen av säkerheten .
koch har producerat ett bra betänkande , emedan det inte har kommit ut mycket av arbetet på cen eller inom ramen för förenta nationernas ekonomiska kommission för europa .
jag vill fråga vice ordföranden om hon i dag kan säga oss hur läget är när det gäller standardiseringssträvandena i dessa båda organisationer samt om eu har möjlighet att snabba på standardiseringssträvandena enligt enklast möjliga principer .
för det står klart att även om vi inför fantastiska bestämmelser här inom europeiska unionen så gör trafiken inte halt vid dessa gränser , den överskrider dem .
därför är det säkerligen meningsfullt med mer långtgående , nämligen regionalt sett mer långtgående regleringar .
om det inte är möjligt att svara på detta i dag , vore det då möjligt att utskottet får ett skriftligt meddelande om hur läget ser ut och hur det står till med förhandlingarna mellan cen och fn : s ekonomiska kommission för europa ?
herr talman ! jag upprepar mina gratulationer till herr koch för hans arbete med det här betänkandet , som på sätt och vis har blivit ett komplement till den debatt vi höll i oktober månad om transport per järnväg .
alla beklagar vi att europeiska standardiseringskommittén ( cen ) inte har haft förmåga att inom de uppställda tidsramarna slutföra den ändring av de bestämmelser som krävs för en lämplig harmonisering inom europeiska unionen .
den här debatten och ändringen av det nu gällande direktivet gör att vi kan ta med andra fakta som visar på mångfalden i vårt europa .
för en stund sedan talade vatanen om låga temperaturer , inte bara om 20 minusgrader utan om 40 minusgrader .
naturligtvis godkänner vi det ändringsförslaget , han har helt rätt , och jag anser att man bör ta med konkreta omständigheter som visar på det varierade klimatet i europeiska unionen , som i vissa fall omvandlas till specificeranden och konkreta krav när man tittar på standardiseringar och karakteriseringar av teknisk art .
vad beträffar swobodas uttalanden om cen : s verksamhet , kan jag tala om att vi har uppmanat dem att påskynda arbetet så mycket som möjligt , för det skulle vara illa om vi , trots den nya fristen , skulle stå inför samma problem om drygt ett år på grund av att arbetet inte har slutförts .
slutligen , herr talman , kan sägas att vi har lyft fram de grundläggande problem som rättfärdigar en ändring av direktivet , vi har talat om förseningen från cen : s sida , om ändringar av vissa bestämmelser , om sambandet mellan direktivets text och innehållet i bilagorna , om behovet av en närmare precisering .
alla bidrag från parlamentets utskott och föredraganden koch , som har omvandlats till olika ändringsförslag , närmare bestämt i fyra , har antagits av kommissionen .
vi godkänner således de fyra ändringsförslag som har lagts fram för oss .
samordning strukturfonderna / sammanhållningsfonden
nästa punkt på föredragningslistan är betänkande ( a5-0108 / 1999 ) av schroedter för utskottet för regionalpolitik , transport och turism om meddelandet från kommissionen om samordning av strukturfonderna och sammanhållningsfonden - riktlinjer för programmen för perioden 2000-2006 &#91; kom ( 1999 ) 344 - c5-0122 / 1999 - 1999 / 2127 ( cos ) &#93; .
herr talman ! det är särskilt tillfredsställande för mig att hålla mitt första tal i europaparlamentet om vad som anses vara den viktigaste frågan i den del av förenade kungariket som jag företräder i detta parlament , dvs. wales .
huvuddelen av wales har , som ni känner till , erkänts mål 1-status enligt strukturfondsprogrammen .
det är helt klart så att många i wales förlitar sig på europeiska unionens strukturfondsprogram när det gäller att lindra en del av de enorma svårigheter som vi utan tvekan står inför .
vi har sett att fattigdomen ökar i wales ; och har ökat ytterligare sedan 1997 .
vi har sett klyftan mellan rika och fattiga vidgas .
vi förlitar oss därför på strukturfondsprogrammen , inte bara för att få till stånd en industriell omstrukturering , utan också för att få till stånd en bredare förbättring av hela den ekonomiska basen i wales .
vad som emellertid är djupt skadligt för oss , är tron att beviljandet av medel från strukturfonderna är något som , på sätt och vis , varit en framgång för regeringen .
det är tråkigt nog bara ett erkännande av de mycket stora svårigheter som wales står inför .
detta är skälet till varför jag vill betona vissa av de frågor som jag anser att kommissionen måste prioritera .
vi vänder oss till kommissionen för att ta itu med frågor som har att göra med kompletterande medel .
vi är missnöjda med det faktum att dessa siffror på något sätt verkar har gömts i förenade kungarikets siffror .
vi vänder oss också till kommissionen för att se till att det finns matchande finansiering för projekten .
vi vänder oss till den för att utmana den brittiska regeringen , för att se till att privata sektorn - som antagligen måste stå för den största delen av utgifterna inom strukturfonderna - deltar vid planeringsstadiet .
vi uppmanar , till sist , kommissionen att se till att pengar från strukturfonderna används på ett öppet och väl redovisat sätt .
alltför mycket av vad som sker i detta parlament är inte öppet och väl redovisat .
detta är ett område inom vilket kommissionen kan hjälpa wales på ett avgörande sätt .
herr talman ! vårt utskott studerar dessa frågor ur många olika synvinklar , men först skall jag tala om forskningens synvinkel .
vi ser mycket positivt på att föredraganden i sina egna slutsatser inkluderat vårt utskotts förslag om att man borde utvidga forskningsinfrastrukturen i sammanhållningsländerna genom att placera ut högskolor och läroanstalter så att de bättre tjänar invånarna i mindre utvecklade regioner och gör det lättare för utbildade personer att stanna kvar i sin hembygd .
detta kan ske genom myndighetsåtgärder , och en sådan decentralisering av den högre utbildningen är utan tvivel nyttig för att utjämna utvecklingen .
en annan fråga som vi uttryckligen skulle vilja belysa ur en industripolitisk synvinkel är att vi gärna sett att kommissionen fäst större uppmärksamhet vid effekterna av ökad användning av tjänster , elektronisk handel och internet när den planerade samordningen av strukturfonderna och sammanhållningsfonden .
tidigare fanns det ett större samband mellan fattigdom / rikedom och näringsstrukturen .
rika var de områden där det fanns arbetstillfällen inom industrin , men i dag har dessa områden kanske blivit till en belastning och kan vara fattiga , vilket gör att man också måste satsa på nya verksamhetsgrenar , på så kallad elektronisk produktion och tjänsteproduktion , eftersom detta är framtidens verksamhetsgrenar .
det ansvariga utskottet har enligt min mening inte i tillräcklig utsträckning tagit hänsyn till detta i sitt betänkande , varför jag å utskottets för industrifrågor vägnar önskar rikta kommissionens uppmärksamhet på denna fråga .
till slut skulle vi i egenskap av utskott för energi ha önskat att man i ännu högre grad framhållit stödet för förnybara energikällor från sammanhållningsfonden och regionala utvecklingsfonden , och därigenom hade man med hjälp av samordning kunnat öka användningen av förnybara energikällor så att energiprogrammets otillräckliga finansiering kompenserats med dessa mer omfattande penningresurser .
( en ) herr talman ! jag vill verkligen tacka fru schroedter för det arbete hon lagt ned i detta sammanhang och förklara för mina kolleger att uttalar mig på min kollega flautres vägnar , som följde detta för utskottet för sysselsättning och socialfrågor , men som tyvärr blivit sjuk .
jag vill rikta uppmärksamheten på ändringsförslag 1 och 2 , vilka röstades igenom av utskottet för sysselsättning och socialfrågor , men inte godtogs av utskottet för regionalpolitik , transport och turism .
dessa ändringsförslag behandlar den sociala ekonomin och behovet av att tillhandahålla socialt riskkapital och finansiellt stödja lokala program för utveckling av sysselsättningsmöjligheter och stärkande av den sociala sammanhållningen .
under årens lopp har parlamentet sett den sociala ekonomin som en viktig och möjlig skapare av arbetstillfällen .
dessa ändringsförslag överensstämmer också med parlamentets syn att social utslagning är en viktig fråga som kräver konstruktiva åtgärder .
vi hoppas att de som överväger att förkasta dessa ändringsförslag har mycket kraftfulla skäl att erbjuda både parlamentet och de medborgare som letar efter arbete .
i sitt betänkande pekade också flautre på ett område inom vilket det i högsta grad saknas samordning , fast detta sannerligen behövs .
i kommissionens förslag hänvisar man till sysselsättningsstrategins fyra pelare och europeiska socialfondens fem åtgärdsområden .
men det är särskilt beklagligt att det här saknas specifika riktlinjer , då idén med att sammanlänka hjälp från socialfonden till sysselsättningsstrategin kommer att träda i kraft för första gången under programperioden 2000-2006 .
man kan säga att denna försummelse ger intrycket att också kommissionen inte har någon idé om hur den skall skapa högsta möjliga samordning mellan hjälp från socialfonden , vilken skall granskas efter tre och ett halvt år , och medlemsstaternas årliga nationella sysselsättningsplaner .
vi hoppas att kommissionen kan ge oss lugnande besked om att detta var ett förbiseende som man nu skall ta itu med på ett konstruktivt sätt .
herr talman , herr kommissionär , ärade parlamentsledamöter ! det förslag som kommissionen har lagt fram av , och därmed uppfyller sitt mandat , betraktar utskottet för jordbruk och landsbygdens utveckling som en vettig utgångspunkt .
men jag vill här poängtera att denna utgångspunkt visar vilka utmaningar vi nu står inför : att förmå befolkningen att stanna kvar på landsbygden , med de förändringar som håller på att ske inom all ekonomisk verksamhet på grund av jordbrukssektorns allt minskande betydelse som inkomstkälla på landsbygden .
detta , tillsammans med bristerna i infrastrukturnätet och samhällsservicen , och arbetstillfällena som i regel är få , ofta säsongsbetonade och tämligen likriktade , ökar flykten från landsbygden .
följderna låter inte vänta på sig .
det är ungdomarna som försvinner , som utbildar sig och får arbete i städerna , något som påverkar landsbygden på ett negativt sätt .
denna bristande infrastruktur är också ett hinder för utbredningen av företag och skapandet av nya arbetstillfällen .
man bör komma ihåg att landsbygden utgör nästan fyra femtedelar av europeiska unionens yta .
inom jordbruket finns endast 5,5 procent av alla arbetstillfällen i unionen .
dessutom driver tre fjärdedelar av alla jordbrukare jordbruk som en deltidssysselsättning och är beroende av ett effektivt tillägg till sina inkomster .
ett av de främsta och viktigaste målen som vi bör fastställa i europeiska unionen är därför att bemöda oss om att skapa nya arbetstillfällen på landsbygden , utanför jordbrukssektorn , inom sektorer som landsbygdsturism , sport , kultur , återerövrande av fädernearvet , omvandling av företag , nya tekniker , tjänstesektorn , etc. även om jordbruket inte längre har en exklusiv roll fortsätter det att vara viktigt , inte bara för att undvika att landsbygden hamnar utanför i ekonomiskt och socialt avseende och att nya spökstäder uppkommer , utan även för att jordbrukarna har en viktig roll i förvaltningen av territoriet , bevarandet av den biologiska mångfalden och skyddet av miljön .
därför förespråkar vi att man fastslår en politik för jordbruket och landsbygdens utveckling som överensstämmer med de mål som vi har satt upp och att landsbygden , i början av 2000-talet , skall vara konkurrenskraftig och mångfunktionell , såväl ur jordbrukssynpunkt som beträffande en öppen attityd gentemot olika verksamheter utanför jordbruket .
det är viktigt att prioritera de allmänna kriterierna för en översiktsplan och befolkningsspridning , och beakta slutsatserna från utskottet för jordbruk och landsbygdens utveckling i fem viktiga avseenden , som endast i viss utsträckning har anammats av utskottet för regionalpolitik , transport och turism under punkterna 16 och 17 .
slutligen vill jag be kommissionen att dessa fem punkter beaktas vid fastställandet av slutsatserna för de fyra pelarna , för jag anser att bevarandet av befolkningen på landsbygden bör vara ett av europeiska unionens främsta mål .
herr talman , herr kommissionär , ärade kolleger ! jag vill börja mitt anförande med att tacka föredragande schroedter för hennes insats .
jag anser att det är ett väl genomarbetat betänkande .
dessutom vill jag tacka henne för hennes vilja till dialog med de övriga politiska grupperna när det var dags att uppnå en avtalslösning inför denna våg av ändringsförslag , som kanske var fler än man hade räknat med , men dessa speglar i själva verket vikten av det betänkande som vi nu diskuterar .
för oss är det viktigt att de slutsatser som antas av parlamentet beaktas av kommissionen , åtminstone andemeningen av dessa , för annars kan det i den här situation verka som att det vi ägnar oss åt är meningslöst och endast en övning i retorik .
faktum är att vi anser , och det framgår av ordalydelsen i slutsatserna , att kommissionen bör ta hänsyn till det som beslutas här i parlamentet , i första hand om granskningen av dessa riktlinjer när halva tiden har gått .
i våra ändringsförslag har vi fastslagit hur viktigt det är att man skapar den nödvändiga samordningen mellan strukturfonderna , sammanhållningsfonden och gemenskapsinitiativen , så att tillämpandet av dessa på bästa sätt , på det mest lönsamma sättet speglar sig i ett successivt utplånande av olikheterna mellan regionerna och i skapandet av sysselsättning , utan tvekan de två viktigaste målsättningarna för de fonder vi talar om .
och som ett sätt att ge en snabb och effektiv impuls till att uppnå dessa målsättningar , anser vi att det är viktigt att de som skapar sysselsättning medverkar i detta initiativ , de som verkligen är driftiga och de som verkligen kan garantera nya arbetstillfällen , det vill säga företagarna .
utdelningen av dessa fonder måste i synnerhet komma de mindre och mellanstora företagen till godo .
om det inte skulle vara fallet , om företagarna känner sig utstötta , om inte företagarna får ta del , och då menar jag inte bara i förvaltningen , utan även i mottagandet av dessa fondmedel , då har vi missat en möjlighet att uppnå våra mål på snabbast tänkbara sätt .
dessutom är det viktigt att vi för att uppnå dessa , för att övervinna olikheterna mellan regionerna och finna källor till sysselsättning , satsar rejält på de nya teknikerna , på näten för transport och kommunikation och på förnybara energikällor .
och detta - jag upprepar - med medverkan av de privata företagen som genom att förena sina insatser med insatserna från den offentliga förvaltningen , som ett komplement till denna utan att det ena för den skull skall hindra eller utesluta det andra , är de som kommer att skapa ett rikt samhälle och nya arbetstillfällen .
herr talman ! det åligger mig att påminna min kollega , evans , om varför wales egentligen erhöll mål 1-status .
det berodde på den skamliga politik som hans eget parti , de konservativa , förde .
låt mig också påminna honom om att när hans partiledare , hague , var wales utrikesminister , bröt han mot varenda regel rörande kompletterande medel , vilket resulterade i ett skarpt formulerat brev från kommissionsledamot wulf-mathies angående föreskrifterna .
jag kan försäkra er om att den brittiska regeringen känner till sina föreskrifter rörande kompletterande medel för mål 1 .
jag föreslår att evans läser bestämmelserna .
min grupp har lagt fram omfattande ändringsförslag till båda de betänkanden som debatteras i dag .
jag vill att vi koncentrerar oss på riktlinjernas avgörande roll .
målet är att tillhandahålla en ram - ett instrument - för stöd och förstärkning av den ekonomiska förnyelsen , för att på ett effektivt sätt använda resurserna i de mest långtgående partnerskapen och att få dessa regioner på rätt köl , så att de kan återhämta sig och få en hållbar utveckling och slutligen kopplas bort från den regionala livsuppehållande apparaten .
det är viktigt att fastställa de kunskaper och möjligheter som finns i våra regioner inom den högteknologiska sektorn .
det är särskilt viktigt mot bakgrund av rapporterna i media som säger att europa snabbt håller på att tappa mark till förenta staterna i de framtida högteknologiska tillväxtbranscherna .
verksamheten inom den förra programrundan visar också på ett tydligt sätt vad riktlinjer inte skall handla om .
de skall inte handla om att skapa ytterligare byråkrati och snåriga bestämmelser .
de skall inte handla om att ändra inriktning och politik när man kommit halvvägs genom projektet , vilket resulterar i oundvikliga förseningar och outnyttjade medel , i synnerhet mot bakgrund av det nya budgetkravet .
tillämpningen och genomförandet av riktlinjerna kan inte överlåtas till personlig tolkning av någon tjänsteman vid kommissionen eller den nationella statliga förvaltningen .
det måste råda en intern sammanhållning vid kommissionsdirektoratet , samtidigt som man respekterar de specifika lokala och regionala aspekterna av kommissionens program .
slutsatsen blir att vi måste se till att riktlinjerna blir breda , vägledande och flexibla för att hjälpa våra programansvariga och de som tar emot medel , och att erhålla maximala möjligheter från våra nya förnyelseområden .
om vi kan tillföra en anda av entreprenörskap i våra fattiga och strukturellt svaga regioner , kommer vi till sist att få dem på rätt köl när det gäller att dra till sig större volymer investeringskapital , som kommer att vara nyckeln till framgång .
det är så vi skall bedöma hur framgångsrika dessa riktlinjer blir : om eu : s regionalpolitik med bra , gedigna och kreativa riktlinjer kan skapa nya möjligheter och göra det möjligt för våra fattiga och strukturellt svaga regioner att efter förmåga bidra till eu : s framtida tillväxt och välstånd .
herr talman , herr kommissionär , bästa kolleger ! jag vill tacka schroedter för ett bra betänkande .
hon har med omsorg satt sig in i ärendet och under utskottsbehandlingen på ett bra sätt beaktat de många ändringar som gjorts i detta betänkande .
föredraganden har också helt riktigt konstaterat att parlamentet inte i tid hörts angående riktlinjerna .
nu är man mycket försenad i frågan .
förhoppningsvis hjälper dock parlamentets ställningstaganden till vid bedömningen av programmen efter halva vägen och vid det praktiska genomförandet av dem .
med tanke på tidpunkten har betänkandet under behandlingen blivit alltför omfattande .
man har där samlat detaljerade frågor och till och med sådant som redan tagits upp i tidigare betänkanden .
i detta skede är det viktigare att koncentrera sig på att bedöma på vilket sätt man genom den här processen skulle kunna styra unionens regionalpolitik med tanke på att målet är att minska den regionala obalansen .
vår grupp framhåller subsidiaritetsprincipen , medlemsstaternas ansvar och de lokala aktörernas roll vid utarbetandet och genomförandet av programmen .
det är speciellt viktigt att involvera de små och medelstora företagen i planeringen och genomförandet av programmen .
vår grupp anser det också vara viktigt att ta mer hänsyn till utomeuropeiska områden och andra ytterområden och vi vill öka växelverkan mellan städerna och landsbygden .
vi motsätter oss ett alltför långtgående förmyndarskap från unionens och medlemsstaternas centralförvaltningars sida och kräver att den byråkrati som fått fotfäste vid utarbetandet och genomförandet av programmen bantas ned .
effekten av projekt som genomförts med hjälp av unionens bidrag har alltför ofta försvagats på grund av långsamt beslutsfattande och krånglig förvaltning .
ofta har man beviljat anslag till projekt som inte gett regionen någon bestående nytta .
projekten måste bli effektivare , mer flexibla och de måste leda till bättre resultat .
i samband med utarbetandet av betänkandet fördes det också en intressant debatt om unionens regionalpolitik i största allmänhet .
det var första gången för oss nya ledamöter och detta är en mycket intressant process .
detta är ett bra betänkande , vår grupp ställer sig bakom det .
herr talman , herr kommissionär , ärade ledamöter ! som ett bevis på att detta parlament ännu inte har kommit över sin roll som rådgivande och underordnad institution , är det utmärkta betänkandet från min gruppkollega elisabeth schroedter ännu inte framlagt i kammaren på grund av att planerna för den regionala utvecklingen under tiden 2000-2006 för mål 1-områden redan har legat flera månader på kommissionens sekretariat .
med hänsyn till detta måste detta parlament hur som helst , innan det godkänner gemenskapens stödramar för den period det gäller , kräva att dessa analyseras och debatteras i kammaren i ljuset av just de inriktningar vi lägger fram i dag , där vi särskilt trycker på deras förmåga att skapa sysselsättning i de fattigaste eller minst utvecklade områdena , och att vi därigenom bidrar till att förändra de nuvarande negativa tendenserna till ojämlikhet i det europeiska samhället och arbetar för ett rättvisare europa .
herr talman ! vi får inte glömma bort att det främsta strategiska målet med strukturfonderna och sammanhållningsfonden och samordningen av dessa är att uppnå en ekonomisk och social sammanhållning .
vi är skyldiga att medverka till utformandet av riktlinjerna och även i utvärderingen av resultaten .
och detta för att vi är medborgarnas företrädare i medborgarnas europa , och inte bara i ett staternas och regionernas europa .
vi kan konstatera att fonderna är en nödvändig , men otillräcklig förutsättning för att uppnå ekonomisk och social sammanhållning .
om vi använder oss av bruttonationalprodukten per invånare som den enda indikatorn kan vi missta oss .
några av kollegerna har redan talat om arbetslösheten , om nedgången i demografin .
vi borde undersöka ett antal indikatorer som tillåter oss att bedöma situationen och utvecklingen i sådana regionala samhällen där situationen är värre än i de övriga .
av vissa av de betänkanden som i dag har lagts fram inför parlamentets plenum framgår det att arbetslösheten i de 25 mest framgångsrika europeiska regionerna är fem gånger lägre än i de 25 minst framgångsrika regionerna .
det tvingar europaparlamentet , herr kommissionären och kommissionen att agera på ett beslutsamt och strategiskt sätt .
jag håller med om att europaparlamentet inte hade någon möjlighet - eller inte fick någon sådan för att mandatperioden snart skulle vara över - att diskutera dessa riktlinjer .
men jag tror inte att betänkandet kommer att dröja .
vi behöver tillsammans fundera över hur de nya programmen med mål 1 och de planer för regional utveckling som har utvecklats innan riktlinjerna träder i kraft , skall kunna bli föremål för en granskning och en riktig utvärdering .
det krävs en samordning av programmen med de olika målen . vi ställer alla kravet att även parlamentet , när halva verksamhetstiden för programmen har gått och det är dags att utvärdera riktlinjerna , skall inta en ledande roll , för vi är medborgarnas företrädare .
medborgarna kan inte acceptera att europeiska unionen fattar beslut på ett så till synes byråkratiskt sätt .
de förväntar sig att den politiska dimensionen finns med , att man visar ansvar , att det finns en kommunikation med medborgarna .
det är det vi i dag vill be herr kommissionären om .
jag hoppas att han , efter sina senaste erfarenheter som regional ordförande , kommer att gå med på att föreslå vissa indikatorer och en strategi till förmån för den ekonomiska och sociala sammanhållningen och inte bara för produktiviteten .
herr talman ! jag stöder huvudförslagen i betänkandet rörande förvaltningen av strukturfonderna och sammanhållningsfonden för perioden 2000-2006 och betänkandets huvudrekommendationer vilka inkluderar följande : det måste alltid råda ett samordnat förhållningssätt till finansieringen ur eu : s strukturfonder och sammanhållningsfonden .
detta innebär att det måste råda ett heltäckande partnerskap mellan lokala myndigheter och nationella regeringar med hänsyn till hur dessa medel skall användas .
medlemsstaterna uppmanas att lägga större vikt vid samordnade strategier för en förnyelse av förhållandena mellan städer och landsbygd .
denna senare fråga är av särskild betydelse .
samtidigt som förnyelsen av våra stadsområden är mycket viktig måste vi alltid hitta en balans i vår politik mellan främjandet av landsbygdens utveckling och förbättringen av livskvaliteten för dem som bor i städerna .
vi har inte för avsikt att bygga ett europa som bara består av städer .
strukturfonderna har spelat en viktig roll för utvecklingen av både städer och landsbygd i perifera länder , huvudsakligen genom förbättring av vägar , vattenrening och transportnät som har samband med detta .
denna process kommer att fortsätta i överensstämmelse med riktlinjerna för finansiella utgifter , vilka fastställdes av eu : s politiska ledare vid toppmötet i berlin förra året , och vilka stöddes av parlamentet vid dess sammanträdesperiod i maj .
tongivande eu-program mellan 1989 , 1993 , 1994 och 1999 har verkligen hjälpt till att förbättra den ekonomiska konkurrenskraften i perifera länder och mål 1-regioner i europeiska unionen .
det viktiga är nu att konsolidera och befästa de framsteg som gjorts hittills .
detta kommer att garantera att randområdena och de yttersta randområdena , de fattigare regionerna i europeiska unionen , hamnar i en ställning där de kan nå framgångar inom det nya euroområdet , såväl som inom den ständigt expanderande inre marknaden där det råder fri rörlighet för varor , personer , tjänster och kapital .
sammanfattningsvis - medan viktiga infrastrukturprojekt fått medel från europeiska regionala utvecklingsfonden och sammanhållningsfonden , bör vi komma ihåg att europeiska socialfonden har spelat en mycket viktig roll vad gäller hjälp till de fattiga i samhället .
socialfonden har verkligen förbättrat våra institutioner för högre utbildning , finansierat våra studieprogram för personer som redan innehar examensbevis och fått till stånd omfattande program som syftar till att bekämpa ungdoms- och långtidsarbetslöshet , hjälpa personer som lämnat skolan vid ett tidigt skede och främja en högre standard vad gäller läskunnigheten hos vuxna .
jag har tidigare flera gånger varit oense med föredraganden , när det gäller regionalpolitiska frågor , men denna gång delar jag hennes uppfattning .
jag vet inte om detta uppmuntrar henne att fortsätta i samma riktning , men i vilket fall som helst skulle jag vilja framföra mina gratulationer .
den andra punkten som jag skulle vilja ta upp är det önskemål som mccarthy och jag framförde i egenskap av föredraganden för den allmänna förordningen . jag skulle alltså föredra att riktlinjerna fogades till förordningen som bilaga .
detta har tyvärr inte skett , och den som bär ansvaret för detta är inte bernié utan det förutvarande utskottet .
jag framför detta för att upprepa parlamentets ståndpunkt .
den tredje punkten som jag skulle vilja ta upp är att jag stöder riktlinjerna i stora drag , i den mån de inte avviker från de anmärkningar vi gjort .
riktlinjerna är till stor hjälp för medlemsstaterna , jag vill särskilt framhålla hur stor betydelse kommissionen tillmäter frågan om hållbar utveckling och ökad sysselsättning , i synnerhet när det gäller likvärdiga möjligheter och transportfrågor .
detta kan åtminstone jag personligen helt och hållet instämma i .
sedan skulle jag i egenskap av öbo vilja kritisera att man försummat frågan om öarnas utveckling .
man lägger inte tillräckligt stor vikt vid detta , och det är heller inte första gången .
under mina fem år som ledamot av parlamentet har jag upprepade gånger berört denna fråga .
herr kommissionär , jag kommer även i fortsättningen att ta upp denna fråga , för i artikel 158.1 i amsterdamfördraget finns en bestämmelse som handlar om en helhetspolitik för öarna .
följaktligen borde kommissionen nu äntligen ta och granska den konkreta frågan .
sedan , herr kommissionär , är det nu äntligen dags att genomföra programmen , även medlemsstaterna måste alltså ta sitt ansvar och sköta sina uppgifter på ett riktigt sätt .
beträffande oss här i parlamentet vill jag påminna om att det finns en uppförandekod för relationerna mellan parlamentet och kommissionen , som undertecknades i maj .
jag är förvissad om att denna kod kommer att följas och att parlamentet kommer att hållas underrättat om detaljer i fråga om genomförandet av programmen .
herr talman ! prioriteringen av ekonomiska kriterier och monetära kriterier ökar orättvisorna i alla dess former .
för den franska planens experter exempelvis är det mest troliga scenariot i dag att de regionala skillnaderna ökar i varje land .
men strukturfonderna har bidragit till att bromsa denna process .
vårt projekt med ett europa som kan uppfylla sociala behov syftar till att höja levnadsstandarden och göra den enhetlig .
genomförandet skulle sannolikt leda till att sådana fördelningsinstrument som strukturfonderna skulle utvidgas .
vi föreslår framför allt en enhetlig kapitalskatt , som skulle göra det möjligt att bidra till fonder som kan åtfölja harmoniseringen av socialförsäkringssystemen och en minskning av arbetstiden på europeisk nivå .
men när kommissionen ombeds att lägga fram riktlinjer gör den det med ett beklagande och på ett luddigt sätt .
det betänkande som i dag läggs fram ger på nytt politiken en plats .
det är ett steg på väg mot en hållbar politik för sysselsättning och utveckling .
och det är det som gör att vi kan rösta för den .
herr talman ! även jag vill tacka föredraganden för ett utmärkt arbete .
mer än någonsin tidigare kommer europa under de kommande åren , på grund av den utmaning som globaliseringen och östutvidgningen medför , att behöva klara och tydliga riktlinjer när det gäller program för att åter få fart på den ekonomiska utvecklingen .
i det avseendet måste europa som helhet , och varje enskild medlemsstat , på bästa sätt utnyttja alla sina resurser och möjligheter , och därmed också de strukturfonder som är tillgängliga .
för att göra det krävs en europeisk kommission som , utöver de goda avsikterna , är tydligare i sina riktlinjer och anstränger sig maximalt i arbetet att kontrollera hur medlemsstaterna utnyttjar dessa resurser .
italien till exempel har under de senaste åren haft problem när det gällt att utnyttja strukturfonderna , framför allt på grund av en överdriven byråkrati , bristfällig information och ett bristande engagemang från de ekonomiska och sociala operatörerna på lokal nivå .
det är därför i första hand två punkter jag vill rikta kommissionens uppmärksamhet på : för det första gäller det att på bästa sätt utnyttja samråd som en metod att samordna lokala och regionala operatörer och göra dem delaktiga i besluten , just för att undvika obalanser och orättvisor .
för det andra måste de administrativa processerna förenklas och göras mer lättillgängliga , eftersom de alltför ofta blir onödigt långa och komplexa , till den grad att de äventyrar tillgången till fonderna , något som framför allt de små och medelstora europeiska företagen klagar över .
herr talman ! låt mig avslutningsvis säga att det är ganska allvarligt att kommissionen i sitt meddelande bara ägnar bristfällig uppmärksamhet åt de territoriella avtalen och framför allt kampen mot arbetslösheten vad gäller kvinnor och ungdomar .
herr talman ! i likhet med min kollega evans , tycker jag att det är synnerligen trevligt att stiga upp i talarstolen och hålla mitt första tal i denna kammare om denna mycket viktiga fråga , särskilt på grund av att jag företräder en del av förenade kungariket , west midlands , som hittills dragit nytta av i synnerhet finansiering från mål 2 .
men det betänkande som behandlas i kammaren i kväll är ett utmärkt exempel på - om vi inte är väldigt försiktiga - hur vi kan lägga fram mycket storslagna idéer som saknar det innehåll som gör dem relevanta för de personer som direkt drar nytta av dem .
betänkandet i sig självt har ett gott syfte men , som så ofta när vi behandlar dessa frågor , saknar ett tydligt syfte och en sund verksamhetsbas .
detta är skälet till varför jag och min grupp lägger fram tre viktiga ändringsförslag och tillägg till texten - inte för att ta bort något från förslaget , utan för att göra det mer relevant för de som det är avsett att ge vägledning .
låt mig förklara hur vi har tänkt här .
för det första vill vi se till att strukturfonderna och sammanhållningsfonden används på ett lämpligt sätt .
erfarenheten visar , i egenskap av företrädare för skattebetalarna i europeiska unionen , att vi bör - att vi måste - kräva finansiell redlighet och öppenhet i samband med utbetalningarna och kontrollen av dessa pengar . våra ändringsförslag och tillägg har därför att göra med uppfyllandet av vad som är känt som &quot; valuta för pengarna &quot; indikatorer under förfarandet där beviljande av anslag sker .
vi får dessutom alltför ofta se att enorma belopp används inom projekt vars resultat man vet kommer att bli otydliga redan vid början av programperioden .
men halvvägs igenom eller vid slutet av denna period finns det inget effektivt sätt att avsluta projektet på , om det inte visat sig vara framgångsrikt .
i våra tillägg uppmanar vi därför till att man skall skapa bestämmelser om strategier för ett praktiskt genomförbart avslutande , så att vi inte bara kan få den nödvändiga garantin mot fortgående kostnader som ofta skattebetalarna får står för , utan så att vi också kan undvika det väl inövade syndromet som innebär att vi offrar ytterligare pengar på ett hopplöst projekt .
slutligen efterlyser vi en förändring vad gäller den balans och den metod som används vid utbetalningen av medel .
det bör vara ett större deltagande från den privata sektorns sida , vilket kommer att ge realistiska ekonomiska perspektiv vid utarbetandet av finansieringsplanerna .
dessutom måste de finansierade projekten - i stället för att vara småskaliga , intäktsbaserade projekt , vilka är svåra att övervaka - bli mer storskaliga , eftersom de positiva effekterna då blir mer uppenbara .
på så sätt kommer det ofta utbasunerade behovet av öppenhet i samband med användningen av dessa medel att minska , och det kommer också frestelsen att i det längre perspektivet på ett onödigt sätt förlita sig på den lokala skattebasen i områden där projekten genomförs . europaparlamentet kommer sålunda att visa hur allvarligt man ser på behovet av sådana reformer .
om dessa ändringar av betänkandet stöds av kammaren i dag , menar jag att detta kommer att förflytta oss till nästa fas , då vi kan åstadkomma de historiska mål som fonderna syftar till , dvs. att på ett ekonomiskt hållbart sätt hjälpa medborgarna i de eftersatta områdena i europeiska unionen att få en tillfredsställande levnadsstandard ; inte genom att ge allmosor , utan att ge hjälp till självhjälp .
jag uppmanar kammaren att stödja dessa ändringsförslag .
herr talman , herr kommissionär , värderade kolleger ! även jag skulle vilja gratulera föredraganden och tacka henne för hennes stora och seriösa arbetsinsats .
det råder inget tvivel om att europeiska unionens strukturpolitik och sammanhållningspolitik är de viktigaste instrumenten för att skapa förutsättningar för utveckling och för att minska de ekonomiska och sociala klyftorna mellan regionerna .
trots de åtgärder som vidtagits består dessa klyftor , och i synnerhet när det gäller arbetslösheten är de mycket större än man kan acceptera .
för att denna politiks mål skall uppnås i största möjliga utsträckning är det nödvändigt att de politiska insatserna samordnas och att de organiseras med ledning av väl genomtänkta , jag skulle vilja säga intelligenta , riktlinjer .
vi får inte glömma att dessa politiska insatser , när de är effektiva , är synliga också för de europeiska medborgarna , som drar nytta av dem och som ser en direkt förbättring av sin livskvalitet .
vi får inte glömma att man särskilt måste uppmärksamma europeiska unionens avsides belägna regioner och dess öregioner , för deras geografiska läge medför stora hinder för deras ekonomiska och sociala utveckling , såvida inte kommissionen kanske har för avsikt att bygga broar eller tunnlar för att förbinda öarna med det europeiska fastlandet .
avslutningsvis skulle jag vilja framhålla att strukturpolitiken i sin helhet måste bli mera flexibel , så att den anpassas till föränderliga situationer och därigenom bättre kan möta de nya utmaningar och nya möjligheter , som uppstår när vi nu har gått in i ett nytt millennium som vi alla knyter varma förhoppningar till .
herr talman ! schroedters betänkande innehåller utan tvivel ganska många viktiga iakttagelser , och därför vill jag gratulera henne .
jag anser emellertid att vi borde hysa ännu större oro när det gäller gemenskapens regionalpolitik , dess inriktning och effektivitet .
man kan sammanfattningsvis konstatera att den enorma massarbetslösheten långt ifrån att lindras tvärtom förvärras ytterligare genom strukturpolitiken .
jordbruksekonomin och jordbruksregionerna drabbas ohjälpligt av den regionalpolitik som bedrivs , med dramatiska följder för sysselsättningen på landsbygden och för jordbrukarnas levnadsvillkor , framför allt i södra europa .
den regionala obalansen ökar dramatiskt inom medlemsstaterna .
om vi betraktar uppgifterna i den sjätte rapporten , skall vi finna att den regionala obalansen har ökat enormt under de senaste tio åren .
man uppmärksammar nästan inte alls de enorma problemen i unionens öregioner , där bristerna i fråga om infrastruktur , transporter , kommunikationer och energi leder till en ständigt fortgående avfolkning .
ansvaret för detta bärs såväl av unionens regionalpolitik som av dess ekonomiska och sociala politik över huvud taget .
stora delar av europas befolkning fördömer skarpt denna politik som farlig och antifolklig .
de nya riktlinjerna har tyvärr samma inriktning , och det finns ingenting som tyder på att inriktningen kan förändras genom att man tillämpar dessa riktlinjer .
herr talman , kära kolleger ! låt mig säga några korta ord för att betona två punkter , som dessa betänkanden påminner oss om , och som har en strategisk betydelse för det perspektiv vi har på unionen .
den första är den väsentliga och centrala betydelse som vi fortfarande fäster vid den ekonomiska och sociala sammanhållningen .
vi oroar oss också över nyheter om att kommissionens känsla för betydelsen av detta mål avtar .
vi kommer att fortsätta att betrakta unionens ekonomiska och sociala sammanhållning som central .
för det andra håller jag med om de ord vi här har hört från en kollega angående öarna , och jag vill även uppmärksamma regionerna i gemenskapens yttersta randområden .
vi skulle i framtiden vilja se mer djärvhet i hanteringen av regionerna i de yttersta randområdena , som beträffande mitt land när det gäller azorerna och madeira .
jag vill passa på detta tillfälle att fråga om kommissionen skulle kunna redogöra för skälen till att kommissionens rapport om gemenskapens yttersta randområden , som parlamentet har väntat länge på , är försenad ?
herr talman , herr kommissionär ! i utskottet för sysselsättning och socialfrågor var vi eniga om kravet på att det viktigaste och strategiskt korrekta var att stödja strukturfondernas och sammanhållningsfondens insatser för en ökad sysselsättning bland de arbetslösa och för jämlikhet mellan kvinnor och män .
tyvärr har inte det kravet beaktats i schroedters utmärkta betänkande , trots att det finns många bevis - något som vi senare kommer att få se i berends betänkande - på hur dessa fonder på ett fantastiskt sätt stöder de sämst utvecklade regionerna att överbrygga det avstånd som skiljer dem från de mest välutvecklade regionerna i europa .
dessa regioner håller på att expandera , vad bni beträffar .
de håller på att expandera i konkurrenskraft , men inte alla får ta del av den ökade rikedomen , för det är inte sysselsättningen som ökar , och skillnaderna i de olika regionerna beträffande arbetstillfällena kvarstår .
herr kommissionär , läs yttrandet från utskottet för sysselsättning och socialfrågor och prioritera detta , för det är där det stora problemet för medborgarna ligger .
och var strategisk i samband med granskningen och beviljandet av fondmedel , och ta hänsyn till behovet av sysselsättning , för det är definitivt något som strukturfonderna och sammanhållningsfonden kräver .
omröstningen kommer att äga rum i morgon kl.12.00.
den sociala och ekonomiska situationen i unionens regioner
nästa punkt på föredragningslistan är debatten om betänkande ( a5-0107 / 1999 ) av berend för utskottet för regionalpolitik , transport och turism om sjätte periodiska rapporten om den sociala och ekonomiska situationen i europeiska unionens regioner &#91; sek ( 99 ) 0066 - c5-0120 / 99 - 1999 / 2123 ( cos ) &#93; .
herr talman , herr kommissionär , kära kolleger ! denna sjätte periodiska rapport om den sociala och ekonomiska situationen i europeiska unionens regioner innebär ett framsteg i analysen av de regionala uppgifterna och belyser vad som hittills åstadkommits på området , sedan den femte periodiska rapporten kom ut .
jag anser emellertid att påståendet att de europeiska regionerna genomsnittligt ligger på samma utvecklingsnivå utgör en något stympad bild av situationen , och tyvärr är det ofta vad som återges i pressen och i vissa tal .
kommissionens rapport sätter till stor del detta påstående i sitt sammanhang , bl.a. när den tar upp den sociala och ekonomiska situationen för vissa regioner inom unionen som ligger mig särskilt varmt om hjärtat : jag tänker på de utomeuropeiska franska departementen och , rent generellt , de yttersta randområdena .
jag gläds därför åt att utskottet för regionalpolitik antagit ett av mina ändringsförslag som uppmanar kommissionen att avsätta ett eget kapitel i den kommande rapporten om sammanhållningen för de yttersta randområdena , närmare bestämt till att analysera effekten av de åtgärder som inom kort kommer att antas genom tillämpning av den nya artikel 299.2 i amsterdamfördraget .
avslutningsvis förefaller det mig som om den sjätte periodiska rapporten innehåller intressanta argument inför ett verkligt projekt för hållbar och rättvis utveckling av det europeiska territoriet , bl.a. när den sammanfattar betydelsen av förhållandet mellan centraleuropa och de yttersta randområdena .
även om kommissionen fortfarande tvekar att säga det alltför tydligt visar den periodiska rapporten att vi snarast måste främja en utveckling av gemenskapen med flera olika utvecklingscentrum , via unionens strukturpolitik och inom ramen för de åtgärder som inletts genom sek ( det europeiska nationalräkenskapssystemet ) .
herr talman ! europeiska socialdemokratiska partiets grupp i detta parlament ställer sig bakom det betänkande som berend just har lagt fram och vi gratulerar upphovsmannen , både till hans fina slutsatser och till hans flexibilitet som har gjort det möjligt för utskottet att införa ändringsförslag från de olika grupperna .
vi bör ha i åtanke att europeiska unionens totala konkurrenskraft utgör 81 procent av konkurrenskraften i förenta staterna , och att denna siffra endast kan förbättras om den gör det i våra konkurrensdugliga enheter , det vill säga i regionerna , och detta i en tid då den tekniska utvecklingen , internationaliseringen av ekonomin och de problem vi har , utvidgningen och den gemensamma valutan kräver en ökad konkurrenskraft av regionerna , men även av företagen och av den enskilde .
europeiska kommissionens sjätte rapport innehåller värdefulla slutsatser .
jag vill sammanfatta två av dessa , som föredraganden redan har tagit upp , en positiv och en negativ sådan .
den första är att betydande framgångar har uppnåtts vad beträffar den territoriella och sociala sammanhållningen i hela unionens territorium , och att gemenskapens fonder har spelat en viktig , om än ej avgörande roll för att minska de regionala olikheterna .
den negativa slutsatsen är att de omfattande insatserna har lett till bättre resultat i fråga om utjämningen av bni och produktiviteten i de europeiska regionerna än i fråga om sysselsättningen .
därför är det viktigt att den strukturella finansieringen i större utsträckning kopplas till skapandet av arbetstillfällen .
det , herr kommissionär , är det främsta budordet för den kommande perioden .
slutligen vill jag , herr talman , uppmana mina kolleger att anta detta betänkande , och i likhet med andra kolleger ber jag kommissionen beakta slutsatserna i den sjätte periodiska rapporten vid utformningen av programmet för åren 2000-2006 .
herr talman , herr kommissionär , bästa kolleger ! för det första vill jag tacka föredraganden för ett bra arbete och också för att han på ett sakligt sätt beaktat ändringsförslagen under utskottsbehandlingen .
den sjätte periodiska rapporten lägger grunden för en bedömning av hur unionens regionalpolitiska mål uppnåtts .
rapporten visar att tillväxten trots alla ansträngningar är ojämn .
den mycket snabba tillväxten i de centrala delarna av europa fortsätter .
de starkaste centra växer också hela tiden snabbare än det europeiska genomsnittet , medan utvecklingen i många sydeuropeiska och nordliga regioner går betydligt långsammare .
nu behövs en djupgående analys av varför regionalpolitiken inte leder till önskat resultat i alla regioner .
är det byråkratin som är boven eller har man inte i tillräcklig utsträckning tagit hänsyn till skillnaderna mellan regionerna , de långa avstånden , det för kalla eller för varma klimatet , den glesa bebyggelsen och de karga förhållandena ?
på vilket sätt kan unionen möta de utmaningar som den globala utvecklingen medför , så att de svagare utvecklade regionerna kan hänga med i utvecklingen ?
det är också viktigt att utreda hur unionens utvidgning kommer att påverka strukturfonderna och utvecklingen av unionens randområden .
medlemsstaterna måste också komma ihåg sitt eget ansvar .
somliga medlemsstater har brutit mot ökningsprincipen och minskat sina nationella regionala medel när regionalstödet från unionen ökat .
detta har tärt på regionalpolitikens resultat .
i fortsättningen måste man också fundera på att utveckla indikatorer för att åtgärderna skall kunna riktas in på rätt plats vid rätt tidpunkt .
man har till exempel inte i tillräcklig utsträckning tagit hänsyn till den okontrollerade migrationen .
även i detta sammanhang finns det skäl att framhålla de små och medelstora företagens avgörande roll som skapare av sysselsättning och som den regionala utvecklingens motor .
alldeles speciellt viktigt är det att överföra den nyaste tekniken och ställa know-how till företagens förfogande i de områden där utvecklingen går långsammare .
vår grupp ställer sig bakom detta betänkande .
herr talman , herr kommissionär , ärade ledamöter ! europeiska unionens regionalpolitik har hittills inte lyckats förändra de befintliga skillnaderna i inkomst per capita .
situationen är allvarlig , vi har alltså i dag i europeiska unionen en tydlig relation mellan arbetslöshet och fattigdom , vilket visas av det mycket oroande faktumet att arbetslösheten uppgår till i genomsnitt 23,7 procent i de mest drabbade regionerna , regioner som sammanfaller med fattiga regioner , medan arbetslösheten i de 25 områden med minst arbetslöshet , vilka ligger i de rika regionerna , bara uppgår till 4 procent .
med hänsyn till denna situation bör behovet av åtgärder ämnade att bekämpa den relativa fattigdomen och arbetslösheten klart framgå i det betänkande parlamentet skall godkänna . åtgärder som exempelvis en riktig tillämpning av strukturfonderna , vilka ofta används felaktigt , för dessa ändamål , genom en central statlig politik , modernisering av telekommunikation och kommunikationer , särskilt genom att integrera de mindre utvecklade områdena i de transeuropeiska järnvägsnäten med inriktning på år 2007 , respekten för och utvecklingen av jordbrukets och fiskets resurser och förmåga i dessa länder , vilka ofta angrips av europeiska unionens egen okänsliga politik , samt främjandet av en aktiv sysselsättningspolitik , framför allt för kvinnor och ungdomar .
bara med en beslutsam tillämpning av denna typ av åtgärder kan man komma över en social och geografisk ojämlikhet som inte är en historisk produkt av oundvikliga misstag , utan tvärtom av en marginalisering och en ekonomisk politik med negativa effekter .
) herr talman , herr kommissionär ! berends betänkande följer exakt den strategi som europeiska kommissionen har definierat genom att frågan om ökad konkurrenskraft ställs i absolut fokus .
det övergripande målet med strukturfonderna , som till exempel skapandet av fler arbetstillfällen , höjd garanti så att alla bereds samma möjligheter , stabilare villkor för sysselsättning och utveckling , nämns endast i förbigående .
detta synsätt förefaller mig oberättigat , och jag ber om att större vikt läggs vid dessa punkter i den sjunde periodiska rapporten .
detta betyder inte att jag inte skulle inse det nödvändiga i att vara konkurrenskraftig , snarare tvärtom i och med att jag själv är företagare i ett mål 1-område , i brandenburg i förbundsrepubliken tyskland , och mycket väl känner till de små och medelstora företagens oro och bekymmer .
i mål 1-regionerna är det parallellt med detta absolut nödvändigt med tidsbestämda åtgärder , och då menar jag åtgärder för att skapa nya jobb , särskilda program för att främja förvärvsarbete bland kvinnor och initiativ för att underlätta för den som vill starta eget .
detta stöds genom lämpliga åtgärder från europeiska unionens strukturfonder .
bara genom att stödja företagens konkurrensduglighet kompenserar man aldrig den eftersträvade sammanhållningen mellan ekonomisk och social utveckling , eftersom det helt enkelt saknas grundförutsättningar för en självbärande utveckling i mål 1-regionerna .
och erfarenheten att den ekonomiska utvecklingen inte själv bidrar till att avskaffa arbetslösheten stöds ju av det faktum att man behöver en ökning av bnp på minst 3 procent för att över huvud taget skapa några nya arbetstillfällen .
den ensidiga koncentrationen på en ekonomisk politik orienterad efter tillgång , efter efterfrågan kan inte fungera så .
och driver man en sådan politik måste man satsa mer på utvidgning och mindre på rationalisering .
man måste absolut länka samman detta med en ekonomisk politik som orienteras efter efterfrågan för att vi alls skall ha en chans att förbättra den sociala situationen i dessa områden .
situationen skiljer sig markant från region till region .
det betyder att det krävs en mängd ytterligare åtgärder för att man alls skall kunna åstadkomma något .
detta vore exempelvis åtgärder för att främja yrkesutbildning , vidareutbildning , för att hjälpa till och slussa tillbaka människor som stötts ut från produktionsprocessen , en flexibel utformning av arbetstid och arbetsformer för att jämka ihop personliga och sociala aspekter på ett avgjort bättre sätt och kanske , återigen , för att främja kvinnors plats i förvärvsarbetet .
herr talman ! mina komplimanger till föredraganden för hans ingående betänkande .
huvudmålsättningen för strukturfonderna är att öka den sociala och ekonomiska sammanhållningen mellan regionerna inom europeiska unionen .
genom att stimulera investeringar av olika slag försöker europeiska unionen att förverkliga en ökning av bnp per capita och en ökning av sysselsättningen .
av den sjätte periodiska rapporten om regionerna kan man dra den försiktiga slutsatsen att dessa stimulanser inte alltid har den önskade effekten .
insatserna som syftar till en ökning av bnp per capita i mål 1-områdena resulterar inte alltid i denna ökning . det kan inte sägas vara ett tillfredsställande resultat under en period där , framför allt under de senaste åren , ekonomisk framgång varit aktuell .
såsom föredraganden anger har dessutom effekterna av strukturåtgärderna varit ringa vad sysselsättningen beträffar .
då är det också på sin plats med en viss återhållsamhet i fråga om gemenskapsstödets effektivitet .
även konstaterandet att skillnaderna mellan regionerna inom medlemsstaterna ibland rentav ökar väcker allvarliga frågor .
herr talman ! det förefaller mig därför vara meningsfullt och nödvändigt att rikta uppmärksamheten , just där det handlar om stimulering av sysselsättningen , såväl på de nationella som på de regionala myndigheterna .
det är ju de som besitter den största kunskapen om de regioner som faller under deras ansvar .
genom att låta dem utveckla skräddarsydda planer för de ifrågavarande regionerna och som komplement till detta , om det är nödvändigt , bevilja ekonomiskt stöd kan man uppnå ett bättre resultat .
och det är ju det som är målet i slutändan .
därför har jag ingenting att invända mot att kommissionen kommer att överlåta det praktiska utarbetandet och genomförandet av åtgärder till medlemsstaterna och regionerna .
det är i anslutning till detta möjligen också mer meningsfullt att över huvud taget lägga en större tyngdpunkt på medlemsstaterna med avseende på det ekonomiska stödet till regioner .
genom att lägga om kriterierna från regionerna till medlemsstaterna förebygger vi en mängd framtida problem .
slutligen vill jag rikta uppmärksamheten på de central- och östeuropeiska ländernas ställning .
av betänkandet framgår det att de i allmänhet ligger rejält efter europeiska unionens länder , i synnerhet på området bnp per capita .
med tanke på den planerande anslutningen inom överskådlig tid för ett stort antal av dessa länder är det absolut nödvändigt att revidera den nuvarande strukturpolitiken .
jag vill härmed , efter andras förebild , också uppmana kommissionen att skyndsamt lägga fram förslag till en revidering .
ärade herr talman , kära kolleger , herr kommissionär ! efter att noggrant ha studerat föreliggande betänkande måste man tvivelsutan dra slutsatsen att det uppsatta målet med strukturpolitiken har kunnat uppfyllas endast till vissa delar .
bland annat har klyftorna mellan regionerna snarare ökat än minskat , medlemsstaterna själva registrerar här ett visst närmande .
likaså har arbetslöshetssiffrorna i de hårdast drabbade regionerna knappast kunnat sänkas , på sina håll har de till och med stigit .
följaktligen frågar jag mig vad det beror på att anslagen från strukturfonderna inte har använts mer effektivt .
inte ens kumuleringen av kapitalet från sammanhållningsfonden och strukturfonderna har varit så framgångsrik i alla regioner som man skulle önska .
eftersom det nu , över hela europa , är alla politikers uttalade mål att sänka arbetslösheten måste man ställa en kritisk fråga huruvida den politik som förs är den rätta eller om det är mindre lämpligt att stärka regionernas konkurrensförmåga genom vederbörliga åtgärder såsom ökat stöd åt forskning och utveckling , förbättrad infrastruktur , höjd utbildningsnivå ?
seriösa strukturreformer och en konkurrensvänligare skatte- och utgiftspolitik är byggstenarna i ett framgångsrikt ekonomiskt säte .
om vi inte vill låta oss förebrås för att driva en kostnadsintensiv strukturpolitik som inte åstadkommer något varaktigt i sysselsättningsfrågan måste vi analysera hittillsvarande åtgärder .
unionens strukturpolitik kan betraktas som framgångsrik i och med att man lyckas skapa tillräckligt många arbetstillfällen och arbetslöshetssiffrorna sjunker markant .
herr talman , herr kommissionär , bästa kolleger ! jag tackar föredraganden för behandlingen av denna mycket viktiga fråga , för den sociala och ekonomiska situationens utveckling kommer att avgöra hur den europeiska allmänheten bedömer att vi har lyckats i vårt arbete .
denna fråga , som påverkar människornas vardag , är en nyckelfråga när det gäller europeiska unionens trovärdighet .
man måste medge att eu redan har stött utvecklingen i fattiga länder , jag skulle till och med säga att den gjort det på ett storslaget sätt .
jag minns hur det såg ut i portugal och i grekland när jag tävlade där för första gången för tjugofem år sedan .
i detta sammanhang säger nog de som talar franska till eu &quot; coup de chapeau &quot; , dvs. jag lyfter på hatten .
eu är verkligen värd en eloge , men skillnaderna mellan fattiga och rika regioner inom länderna är fortfarande för stora .
vad blir konsekvensen ?
folk reagerar genom att rösta med fötterna , genom att ge sig iväg , på jakt efter bröd .
därför tvingas vi att för samma människor i ett och samma land bygga skolor , sjukhus , hela infrastrukturen om och om igen .
detta är oerhört dyrt och skapar också mycket stora sociala problem .
de allra flesta skulle dock vilja bo kvar i sin födelsebygd om de fick möjlighet till det , dvs. om det fanns arbete där .
vi måste ge dem denna möjlighet .
detta är eu : s och vår moraliska skyldighet .
som lösning ser jag en klar uppmuntran till företagsamhet .
med företagsamhet menar jag ingalunda bara att man äger ett företag utan jag menar ett viljemässigt tillstånd .
jag menar den inställningen att en människa vill gå framåt i sitt liv oavsett om hon är arbetare , företagare eller tjänsteman .
hur ser ett rättvist samhälle ut ?
ett samhälle där en människa från enkla förhållanden kan gå framåt i sitt liv för att hennes barn skall få det litet lättare .
på det sättet är det också möjligt att utveckla regionerna i en positiv riktning , för människorna är företagsamma och arbetar om man ger dem möjlighet till det .
avslutningsvis skulle jag vilja säga att vi i detta fall borde ta lärdom av amerika där fliten fortfarande står högt i kurs och framgång är ett bevis på kompetens och inte ett föremål för avundsjuka , som ofta är fallet hos oss i europa .
herr talman , herr kommissionär , kära kolleger ! eftersom jag har begränsat med tid skall jag bara ta upp det viktigaste .
vi kan först och främst konstatera att resultatet av tillväxten inte är rättvist fördelat inom unionen .
ett exempel är de yttersta randområdena , som fortfarande är hårt drabbade av mycket hög arbetslöshet .
la réunion har exempelvis en arbetslöshet på 37 procent .
men det beror inte på konjunkturen utan det är fråga om en strukturmässig arbetslöshet . den skapas av det faktum att vi befinner oss långt bort och är en öregion , kort sagt det beror på vår personlighet .
för att bemöta detta innehöll artikel 299.2 i amsterdamfördraget en princip om särskild och undantagsmässig behandling .
nu återstår att omsätta denna princip i handling .
kommissionens dokument som skulle komma i december 1999 har skjutits upp till januari och sedan till februari , och de första kommentarerna gör mig knappast optimistisk .
jag vänder mig därför högtidligen till rådet och kommissionen .
när det gäller skattefrågor , statligt stöd , strukturfonderna eller att försvara våra traditionella produkter måste vi snarast utarbeta konkreta åtgärder som är både djärva och ambitiösa .
annars kommer konvergens och sammanhållning tyvärr bara att vara tomma ord , och det finns risk för att den strukturpolitik som bedrivs i våra regioner slutar med ett misslyckande trots att det handlar om så stora belopp .
( fr ) herr talman ! jag skulle i min tur , liksom alla andra talare , vilja tacka herr berend och lyckönska honom till ett utmärkt arbete .
liksom när det gäller det tidigare betänkandet är analysen mycket kompetent och exakt , och rekommendationerna , liksom era egna kommentarer mina damer och herrar , kommer att vara till nytta för kommissionen i allmänhet , och för kommissionären med ansvar för regionalpolitik i synnerhet , när vi skall inleda programplaneringen i fråga om anslagen för 2000-2006 .
jag skulle i min tur vilja göra några kommentarer , till att börja med om er bedömning , herr föredragande , av denna sjätte periodiska rapport .
ni betonade dess kvalitet och ni skrev till och med , om jag inte misstar mig , att i jämförelse med de tidigare var den betydligt bättre .
jag vill för kommissionens räkning och för min företrädares , wulf-mathies räkning , säga att vi var mycket glada över denna bedömning från kammaren och er .
kommissionen har verkligen ansträngt sig , herr berend , för att denna sjätte periodiska rapport skulle göra det möjligt att konstatera en insats , ett kvalitativt steg framåt , i den analys vi föreslår er .
jag tänker särskilt på innehållet i kapitel 2.1 i rapporten , där kommissionen på ett fördjupat sätt granskat de ekonomiska definitionerna av den regionala konkurrenskraften och försökt analysera hur denna konkurrenskraft kan stödjas , förbättras och påverkas av faktorer som vissa av er , markov nyss eller raschhofer , kraftigt betonat .
jag tänker på teknisk forskning och utveckling , infrastrukturens tilldelning och kvalitet , de mänskliga resursernas potential , de små och medelstora företagen och direktinvesteringar från utlandet .
så långt kvaliteten .
herr föredragande ! jag vill inte nu lägga alltför mycket tid på detaljer om min uppfattning inom olika allmänna punkter där kammaren redan är överens med oss .
jag skall bara kort nämna dem : den första gäller betydelsen av rapportens slutsatser för att utarbeta prioriteringar för den nya regionalpolitiken , särskilt för förhandlingar om programplaneringsdokument med medlemsstaterna .
den andra punkten , partnerskapen , som flera av er betonat , handlar om rollen för de lokala och regionala myndigheterna , den privata sektorn , arbetsmarknadens parter samt föreningarna och lokala grupper .
när det gäller problemet med partnerskap kommer jag att mycket noggrant se till att bestämmelserna i den allmänna förordningen om strukturfonderna tillämpas korrekt .
den tredje punkten gäller behovet av att öka sysselsättningens andel av tillväxten , även om jag mycket väl vet , och van dam sade det också nyss , att det i första hand är medlemsstaterna som är ansvariga , och att man , när man talar om medlemsstaternas ansvar , liksom om nyttan och effektiviteten av denna regionalpolitik , också måste titta på var vi befinner oss .
fruteau förklarade nyss att resultatet av tillväxten är orättvist fördelat .
herr parlamentsledamot ! det måste ändå finnas en tillväxt och vi kan inte befinna oss i en period av fullständig stagnation eller tillbakagång , vilket förekommit tidigare .
tillväxt och fattigdom gäller inte alla , kanske ni hävdar .
när tillväxt är ett faktum måste den vara bättre fördelad , men det som är ännu svårare och drabbar de regioner som är avlägset belägna , de yttersta randområdena eller öregionerna ännu allvarligare , är avsaknaden av tillväxt som varit kännetecknade för de två senaste decennierna .
den fjärde punkt som hedkvist petersen nyss betonade är främjandet av en politik för lika möjligheter för män och kvinnor .
den femte punkten gäller de små och medelstora företagens betydelse och roll , vilket vatanen starkt betonade nyss .
slutligen har vi den positiva effekten av strukturfondernas förvaltningssystem på de nationella myndigheterna , tjänstemännens motivation när de förvaltar dessa fonder , även om det ibland är komplicerat , och betydelsen av att på nytt förbättra förfarandet för kommissionens utvärdering , uppföljning och kontroll .
jag vill i det sammanhanget informera europaparlamentet om min avsikt att i mitten av år 2000 arrangera ett seminarium med nationella och regionala myndigheter om denna fråga om utvärdering av förfarandena för utbyte av goda tillämpningar när det gäller att förvalta strukturfonderna .
herr berend ! ni ville att zonindelningen skulle genomföras snabbt .
vi har avslutat den .
i morgon kommer fyra nya länder att vara föremål för kommissionens beslut och mycket snabbt , hoppas jag , är det italiens tur .
ni kommer alltså att bli nöjd på den punkten eftersom alla länder som berörs av mål 2 blir indelade i zoner .
när det gäller den informella ekonomin som ni tar upp i ert betänkande , vet jag naturligtvis att analys och framtagning av statistik på detta område är beroende av uppgifternas tillförlitlighet och såsom cocilovo också sade föreligger det ett tillförlitlighetsproblem när det gäller dessa uppgifter .
i viss utsträckning beaktas de på nytt i statistiken över bni och undersökningar om arbetskraften och i vilket fall som helst vill jag betona de ansträngningar eurostat gör och kommer att göra för att förbättra statistikens kvalitet .
herr berend ! liksom aparicio sánchez tog ni upp avsaknaden av reformer på fiskeområdet .
på denna punkt , som personligen intresserar mig , vill jag erinra om att denna sektor är liten - vilket inte betyder att den är betydelselös - och att den är koncentrerad till ett mycket litet antal regioner , och det gör det inte lättare att analysera den inom en regional ram .
denna typ av sektorsanalys faller mer under generaldirektoratet för fiske , under min kollega fischlers ledning .
jag vill ändå försäkra er om att kommissionen kommer att försöka införliva en sådan analys i den andra rapporten om sammanhållningen , som sannolikt bättre kommer att motsvara denna oro .
flera av er har nämnt punkter som bör ingå i denna andra rapport om sammanhållningen , och föredraganden tog upp några av dessa .
jag vill till att börja med försäkra er om att sammanslagningen av de periodiska rapporterna och rapporten om sammanhållningen inte på något sätt kommer att innebära att information går förlorad eller att intresset minskar för innehållet i rapporten om sammanhållning som för mig , herr föredragande , är ett mycket viktigt instrument , inte bara för att man redogör för vad som gjorts och gör det på ett öppet och noggrant sätt , eller för att man granskar eller utvärderar kommande riktlinjer , utan också för att skapa en allmän debatt med medborgarna och även med er som folkvalda om denna regionalpolitik och om det som en dag skulle kunna bli en europeisk politik för fysisk planering .
jag har i vilket fall som helst noterat att ni önskar införliva följande punkter i rapporten : definition , insamling och analys av beståndsdelar som är representativa för regionen och för alla länder i central- och östeuropa , ett kapitel om de yttersta randområdena och öregionerna som flera av er tagit upp , särskilt sudre och fruteau , analys av regionernas konkurrenskraft i länderna i central- och östeuropa - det blir den stora utmaningen för oss , för er , för kommissionen , under de kommande åren , och slutligen de gränsöverskridande aspekterna .
på alla dessa punkter skall jag försöka följa era rekommendationer .
jag skulle slutligen vilja ta upp några politiska slutsatser som ni för övrigt känner till , men där jag ändå skulle vilja erinra om de viktigaste beståndsdelarna .
mina damer och herrar ! avsevärda framsteg har gjorts för att uppnå en verklig konvergens , bl.a. för de fyra sammanhållningsländerna , men också , herr pohjamo , det säger jag ärligt , för regionerna inom mål 2 som tagit igen viss försening i sin utveckling , bl.a. när det gäller infrastruktur .
det är den första politiska punkten .
den andra politiska punkten , strukturfonderna , har lämnat och kommer att lämna ett betydande bidrag till denna tillnärmningsprocess .
alla makroekonomiska modeller som vi arbetar efter visar för det senaste decenniet att mer än en tredjedel av den konvergens som uppnåtts i regioner med försenad utveckling inte skulle ha ägt rum om det inte vore för strukturfonderna .
jag har emellertid noterat , när det gäller framför allt de yttersta randområdena , fru sudre , herr fruteau , och även herr nogueira román , att ni konstaterar att mycket fortfarande återstår att göra - och det är min tredje punkt - när det gäller att öka sysselsättningen , förbättra kampen mot social utslagning , som är särskilt allvarlig och oacceptabel i många av våra regioner samt underlätta för kvinnor och ungdomar att komma in på arbetsmarknaden .
den fjärde politiska punkten gäller unionens utvidgning , som är det stora politiska och humanistiska projektet för våra institutioner under de kommande åren , och även en stor utmaning för europas sammanhållningspolitik , en punkt som van dam betonade .
jag tror att redan i berlin och i de finansiella instrument som ställs till vårt förfogande kan man ana det som skulle kunna bli en sammanhållningspolitik för de första nya länder som skall bli medlemmar .
jag tänker särskilt på ispa-instrumentet som det är mitt ansvar att genomföra under de kommande veckorna .
mina damer och herrar ! som ni ser har vår nya programplanering knappt inletts och vi har redan en gemensam diskussion om effekten av unionens utvidgning på vår strukturpolitik .
denna sjätte periodiska rapport som ni , herr berend , totalt sett uttalat er positivt om utgör för oss , för mig , en bra bas för diskussionerna .
jag skulle därför vilja tacka er mycket uppriktigt för ert bidrag till diskussionerna som vi inlett för de kommande riktlinjerna , liksom för den goda tillämpningen av riktlinjerna för perioden 2000-2006 .
( sammanträdet avslutades kl. 20.25 . )
tack så mycket , herr cox !
jag förstår vad ni menar .
vi har noterat det .
herr talman ! beträffande punkt 11 i arbetsplanen kom vi i går överens om att bourlanges betänkande skulle vara med på dagens föredragningslista .
emellertid drogs det tillbaka av budgetutskottet i går kväll utan att diskuteras eller bli föremål för omröstning .
det måste därför strykas från dagens föredragningslista .
. herr wynn , det är logiskt .
betänkandet har följaktligen avförts från föredragningslistan .
herr talman ! vad beträffar lynnes kommentarer i går om hälsa och säkerhet i denna byggnad antar jag att hon talade om avloppet , för det finns en hemsk kloaklukt på femte våningen i tornet .
detta måste undersökas eftersom det är ett klart tecken på att någonting är väldigt fel .
jag vill inte komma dragande med frågan om denna byggnad i all oändlighet , men detta är ett allvarligt problem .
. fru ahern , vi har noterat det .
jag vill be er att lägga fram detta speciella fall , som rör fläktarna på en viss våning , för kvestorerna , eftersom de egentligen är ansvariga för det .
men vi skall också vidarebefordra det till våra enheter .
reformering av den europeiska konkurrenspolitiken
herr talman , herr kommissionär ! vi för i dag en viktig debatt om europeiska unionens konkurrenspolitik .
vi diskuterar en mycket omstridd modernisering av den europeiska kartellrätten , nämligen wogaus betänkande , och den är mycket mer omstridd än kanske omröstningen i utskottet för ekonomi och valutafrågor gett vid handen .
jag vill absolut säga att jag personligen anser att kommissionens förslag i detta konkreta fall är felaktigt , och att det återstår att se huruvida begreppet modernisering verkligen är befogat för vitbokens innehåll i artiklarna 81 och 82 , eller om inte snarare begreppet tillbakagång vore mer tillämpligt i detta fall .
vi talar i dag emellertid också om översikten över statligt stöd och den allmänna rapporten om konkurrenspolitiken för 1998 , där mitt inlägg i denna gemensamma debatt gäller det senare området .
men båda områdena - rapporten om konkurrenspolitiken och översikten över det statliga stödet - har naturligtvis också en gemensam grundval i denna vitbok .
det gäller kravet på modernisering , på den europeiska konkurrenspolitikens framtidsförmåga .
om man läser kommissionens båda dokument ser man att 1998 var ett år där man fortsatt den modernisering som inletts under 1997 och delvis också avslutat den ; det känner vi själva till från vårt löpande parlamentariska arbete .
låt mig göra två principiella påpekanden : kommissionen har , som ansvarig myndighet , med sin konsekventa hållning alltid gjort stora insatser för konkurrensfriheten , inte alltid till glädje för berörda medlemsstater eller företag .
den bör fortsätta på denna väg .
men , herr kommissionär , allt detta blir i framtiden inte mindre komplicerat - jag vill bara erinra om utmaningarna på grund av utvidgningen av unionen , fördjupningen av den inre marknaden , de tekniska framstegen och globaliseringen .
det hänger faktiskt inte bara på moderniseringen av gemenskapsrätten , utan det beror mer än någonsin på öppenheten i besluten i de enskilda fallen , och på möjligheten att även kunna sätta sig in i besluten , ty den europeiska konkurrenspolitiken kommer att vara beroende av acceptansen från befolkningen , liksom från de berörda politiska instanserna och företagen .
men - utan öppenhet ingen acceptans , och då alltså inte heller någon modernisering utan öppenhet .
rapporten om konkurrenspolitiken 1998 är inte någon dålig grundval för detta , men det finns inte heller någonting som inte skulle kunna göras bättre .
en rad impulser kommer vi att lämna vidare till er , herr kommissionär , tillsammans med vår resolution , men en delaspekt vill jag redan nu gå in på : öppenhet och redovisningsskyldighet hör ihop .
jag vill inte rubba ansvarsfördelningen mellan kommissionen och parlamentet .
kommissionen är det verkställande organet , och parlamentet bör för sitt eget oberoendes skull inte heller vilja vara det , utan parlamentet är ett kontrollorgan , och var kan man bättre klargöra bakgrunden till sina beslut än i det demokratiskt valda parlamentet och just i en ständig parlamentarisk diskussion ?
även här bör vi fortsätta på den inslagna vägen , intensifiera den och göra den beständig .
men en sak vill jag säga helt tydligt : parlamentet är lagstiftande , och att vi just när det gäller konkurrensrätten bara har samrådsrättigheter , är egentligen skandal !
här riktar vi ett krav till rådet och regeringskonferensen att införa ett medbeslutandeförfarande när det gäller konkurrensrätten .
jag förväntar mig av kommissionen att man fullständigt utnyttjar alla möjligheter till parlamentarisk medverkan , om det finns tvivel om att parlamentet skall kunna delta , och detta också redan i den fördragssituation vi har nu .
jag förväntar mig också att kommissionen kommer att stödja oss offensivt i fråga om kravet på medbeslutande i lagstiftningsförfarandet .
det kommer att utgöra ett prov på hur klokt våra institutioner kan samarbeta .
trots att man bekänner sig till konkurrensprincipen är konkurrensen dock inte något mål i sig .
konkurrens är ett instrument och leder inte alltid till optimala lösningar .
det hör nu en gång till de elementära kunskaperna i ekonomi att marknaden i många avseenden misslyckas , och den som bestrider detta är en ideolog , och ingenting annat .
konkurrensen skall balansera utbud och efterfrågan , och sörja för en optimal fördelning av de ekonomiska resurserna .
men en optimal effektivitet inställer sig inte nödvändigtvis av sig själv .
det krävs ramvillkor för att förhindra missbruk , till exempelvis genom kartellrätten .
men därmed förhindras huvudsakligen endast missbruk , det räcker inte ensamt till för att uppnå de mål som legitimeras av samhället .
ja till konkurrens , och en inskränkning av stöden där så krävs och där det är möjligt !
men eftersom stöden i rapporten om konkurrenspolitiken 1998 utgör den största delen vill jag , oaktat kollegan junkers betänkande , ändå tillfoga följande : stöd till små och medelstora företag när det gäller forskning och utveckling , när det gäller utbildning i regionalpolitik och miljöpolitik , det är absolut möjligt och måste också vara genomförbart .
stöd måste tillåtas just för sådana mål , så länge de inte leder till oacceptabla snedvridningar av konkurrensen .
just här är det ännu viktigare att besluten är förståeliga än i fråga om kartell- och fusionsrätten .
stöden bör inte nedvärderas , utan man måste se på hur de kan bidra till att man uppnår de mål som just nämnts .
det sista påpekandet riktade sig mindre till kommissionen , utan snarare till kollegerna i ppe-gruppen .
herr talman , herr kommissionär , mina kära kolleger ! det betänkande som jag i dag har tillfälle att lägga fram för er , är ett yttrande om kommissionens årliga rapport över statliga stöd inom europeiska unionen , för vilka gemenskapen är behörig i kraft av artiklarna 87 , 88 och 89 i fördragen .
kommissionens rapport är i huvudsak beskrivande ; här redogörs för statsstödens utveckling såväl inom tillverkningsindustrin som inom andra sektorer , enligt kriterier som finansieringsmetoder och eftersträvade mål .
när det gäller rapportens kvantitativa avsnitt tillåter jag mig att hänvisa till motiveringen . här nöjer jag mig med att peka på att årsbeloppet i genomsnitt ligger på 95 miljarder euro för perioden i fråga , vilket utgör en minskning på 13 procent i förhållande till perioden 1993-1995 , något som i huvudsak beror på en minskning av stöden i förbundsrepubliken tyskland .
i klartext ligger de anmälda statsstöden i stort sett på ett stabilt genomsnitt under den granskade perioden , och tar ungefär 1,2 procent av gemenskapens bni i anspråk . det motsvarar händelsevis mer eller mindre gemenskapens budget för ett år .
samtidigt är skillnaderna mellan staterna avsevärda och kan bedömas på olika sätt , bl.a. i procent av mervärdet och per löntagare .
det kan också vara av intresse att lägga till de statliga stöd och gemenskapens interventioner som på något sätt kan likställas med statsstöd .
då framgår det klart och tydligt att det är de fyra länder som bl.a. får stöd från sammanhållningsfonden som hamnar i toppen av klassificeringen .
därmed kommer jag fram till betänkandets förslagsdel .
vi kan först och främst konstatera att kommissionen anser att informationen ( såsom den presenteras i kommissionens årliga rapport ) täcker alltför stora områden för att tillåta en grundligare utvärdering av statsstödspolitiken , något som är såväl berättigat som förnuftigt med hänsyn till nationella intressen , och mycket viktigt med avseende på respekten för konkurrensen , enligt definitionen i fördragets bestämmelser .
kommissionen kan endast samla in och analysera de uppgifter som medlemsstaterna anmäler .
det är således staternas och regionernas sak att garantera kvaliteten på de uppgifter som lämnas in , och vårt utskott anser att man bör göra ytterligare insatser för det ändamålet .
av samma skäl försvarar vårt parlamentsutskott det redan gamla förslaget om ett offentligt register över statsstöden , som bl.a. skall finnas tillgängligt på internet .
om uppgifterna blir bättre och mer detaljerade , i synnerhet i förhållande till eftersträvade mål och noterade resultat , kommer europeiska kommissionen själv att kunna företa , eller låta företa , regelbundna studier för en social och ekonomisk utvärdering av nationella och regionala stöd .
i den mån sådana studier redan finns , bör kommissionen så öppet som möjligt informera om dess egna synpunkter i förhållande till fördragens mål , som inte bara är att säkerställa den europeiska ekonomins konkurrenskraft , utan också en hållbar utveckling och ekonomisk och social sammanhållning .
genom att i första hand lägga tonvikt på kvaliteten på den information som lämnas , har vårt utskott undvikit att - i våra debatter och därmed i det betänkande som jag har äran att presentera för er - göra det enkelt för oss genom att i förväg hävda att statsstöden i sig är alltför stora alternativt otillräckliga .
en majoritet av utskottets ledamöter har i stället strävat efter en jämvikt ; å ena sidan bör man kräva att såväl staterna som företagen respekterar konkurrensreglerna och å andra sidan bör man erkänna att den här typen av stöd kan medverka till att fördragets mål förverkligas , i synnerhet , som jag redan har nämnt , i fråga om hållbar utveckling , forskning och utveckling samt ekonomisk och social sammanhållning .
samtidigt har utskottet godkänt en rad olika ändringsförslag till föredragandens ursprungliga utkast , vilka bl.a. betonar att stöd som bedöms vara illegala skall betalas tillbaka och att det upprättas en resultatlista .
sju ändringsförslag har givits in på nytt inför det här plenarsammanträdet .
flertalet av dem förmedlar våra politiska skiljelinjer i fråga om statsstödens lämplighet och effektivitet , med tanke på att enbart privata investeringar inte räcker till , vare sig detta medges eller ej , market failures eller marknadens otillräcklighet .
det finns bl.a. ett ändringsförslag rörande energisektorn , som jag i egenskap av föredragande vill framhålla som särskilt betydelsefullt .
herr kommissionär ! jag vill avsluta denna presentation genom att å ena sidan framhålla ett orosmoln och å andra sidan en begäran från ledamöterna i vårt utskott .
oron avser de central- och östeuropeiska ländernas anslutningsprocess i förhållande till konkurrenspolitik och statsstöd .
detta är med största sannolikhet en komplicerad fråga , och vi skulle önska att kommissionen redogjorde för sakens nuvarande läge , bl.a. vad gäller de ansökande ekonomiernas kapacitet att respektera konkurrensreglerna , och när det gäller statsstöd ; det sannolika behovet av att fastställa specifika regler om statsstöd för en omstrukturering av deras sektorer .
till sist , och härmed skall jag avsluta , en begäran som rör europaparlamentets framtida behörighet inom de områden som vi nu talar om - konkurrenspolitik och statsstöd - en möjlighet med tanke på nästa regeringskonferens .
som ni vet , herr kommissionär , försvarar vi i detta betänkande tanken att medbeslutandeförfarandet skall tillämpas för grundläggande lagstiftning om statliga stöd .
min del i dagens debatt gäller gemenskapsreglerna för stöd till stålindustrin . det är det allmänna stödet som lämnats i europa i enlighet med dessa gemenskapsregler , och som kommissionen har granskat .
det är totalt 27 fall under år 1998 . dessa fall har kommissionen avgett en egen rapport om .
eksg-fördraget kommer att löpa ut inom kort .
den fråga som vi i dag i synnerhet måste ägna oss åt är hur stödet till stålindustrin skall hanteras i framtiden .
kommissionens beslut , som framläggs i översikten , välkomnas av europaparlamentet , inklusive beslutet att i ett konkret fall kräva tillbaka medlen med tillämpning av artikel 88 i eksg-fördraget .
den europeiska stålindustrins konkurrenskraft behandlas samtidigt också i kommissionens senaste meddelande , som vi ännu inte har diskuterat i parlamentet .
liksom på andra områden gäller även för järn- och stålindustrin ett generellt förbud mot stöd enligt artikel 87.1 i eg-fördraget .
enligt denna artikel är statligt stöd principiellt oförenligt med den gemensamma marknaden .
undantag tillåts endast i exakt definierade fall .
enligt artikel 88 är kommissionen ålagd att kontrollera statliga stöd .
år 1998 var det viktigaste fallet när preussag i tyskland försågs med kapital till ett belopp av 540 miljoner euro .
dessutom måste medlemsstaterna meddela kommissionen sina stödåtgärder i förväg .
vad beträffar stålindustrin ställdes de gällande reglerna upp den 18 december 1996 .
enligt dessa kan stöd till förmån för stålindustrin endast lämnas i bestämda , exakt definierade fall . det är forsknings- och utvecklingsstöd , miljöskyddsstöd , socialt stöd vid stängning av stålverksanläggningar och stöd för den slutliga nedläggningen i icke konkurrenskraftiga företag .
dessutom finns det en särbestämmelse om upp till 50 miljoner euro för medlemslandet grekland .
uppenbarligen har det under de gångna åren ändå uppstått problem i den praktiska hanteringen av gemenskapsreglerna till stöd för stålindustrin , som inte har tagits upp fullständigt i betänkandet .
ur parlamentets synvinkel är det viktigt att man redan i dag talar om bestämmelser som kan träda i kraft när dessa gemenskapsregler för stöd till stålindustrin har löpt ut .
det får inte beslutas om någon uppmjukning av befintliga grundvalar för gemenskapsreglerna för stöd till stålindustrin .
ingen vill ha en hämningslös subventionskonkurrens i europa .
detta skulle avsevärt skada den inre marknaden även efter den konsolidering av stålindustrin som skett under de senaste åren .
därför anser parlamentet att det är nödvändigt att bestämmelserna om subventioner till stålindustrin ändras med tanke på skillnad i behandling som industrin påstår har ägt rum , och att kommissionen för rådet lägger fram bestämmelser som skall träda i kraft när de nuvarande bestämmelserna löpt ut .
vi känner till att rådet hittills vägrat besluta om sådana bestämmelser .
det beror också på att man tror att man , när gemenskapens regler om stöd till stålindustrin löper ut , återigen kan göra som man vill , utan den besvärliga kontrollen från kommissionens sida .
vi kräver därför att gemenskapsreglerna om stöd till stålindustrin skall regleras genom en förordning från rådet enligt artikel 94 när fördraget löpt ut , eftersom de endast på så sätt kan bli klara och rättsligt bindande .
det strikta förbudet mot allt stöd , som inte täcks av gemenskapsreglerna , kan bara iakttas på detta sätt .
en förordning från rådet , som omedelbart träder i kraft , måste också iakttas av de regionala regeringarna .
även i framtiden måste vi undvika intrång i konkurrensvillkoren och störningar i balansen på marknaderna .
man måste också kritisera kommissionens praxis att godkänna upprepat stöd för stålföretag , som enligt kommissionens åsikt inte faller under kategorierna i gemenskapsbestämmelserna , även om eg-domstolen i enstaka beslut har godkänt denna skillnad i behandling .
i ett betänkande som återstår att utforma för år 1999 uppmanas kommissionen att detaljerat klarlägga sin aktiva roll vid utarbetandet av omstruktureringsplaner och godkända undantagsfall , och därmed på denna grundval möjliggöra en korrekt utvärdering av de totala sammanhangen .
efter att utskottet för ekonomi och valutafrågor enhälligt har antagit förslaget till betänkande , med två nedlagda röster , ber jag att vi i kammaren helt och fullt godkänner denna framställning , som vi själva har initierat .
herr talman , kära kolleger ! den inre marknaden är inte fullbordad .
subventioner , monopol och konkurrenshinder hämmar fortfarande både marknader och utveckling .
nationella regeringar skjuter till subventioner och lovar att det är sista gången , men så upprepas det igen .
subventioner snedvrider allokeringar , både inom och mellan länder .
en successiv avveckling av statsstödet behövs , och alltfler marknader måste öppnas för konkurrens .
det gäller både dem som har monopoliserats privat och offentligt .
offentliga monopol avvecklas oftast motvilligt .
ökad konkurrens och nyetableringar skulle kunna ge betydande välfärdsvinster - även inom utbildning , sjukvård och social service .
offentliga monopol måste ersättas av konkurrenskraftiga strukturer .
europa måste moderniseras och anpassas till entreprenörskap och en konkurrenskraftigare miljö för konsumenter och företag .
effektiv konkurrens pressar priser och höjer levnadsnivåer .
konsumentpolitiken har i alltför liten utsträckning inriktat sig på just prisnivåerna .
konkurrenspolitik och konsumentpolitik hör ihop .
inre marknaden är grunden för vårt arbete .
dess lagstiftning skall gälla lika för alla , för stora som för små länder .
en systematisk genomgång av de nationella regelverken behövs för att undanröja konkurrenshinder .
även eu : s eget regelverk kan då behöva en analys .
den nya modell som nu prövas av kommissionen får inte leda till en ren nationaliseringsprocess som skulle urholka den uppnådda konkurrenspolitiken .
den måste vara väl förankrad i medlemsstaternas nationella myndigheter för att bli effektiv .
om ett halvår kan det vara lagom att göra en analys av utfallet , men även att se närmare på den nya situationens effekter på kommissionens roll .
tanken på att hålla en institutionellt övergripande kongress som öppnar för en förutsättningslös debatt utifrån ett brett perspektiv med representanter från olika intressenter har tills vidare löst frågan om hur man skall gå vidare .
då finns det tillfälle att slå fast nya principer eller återkomma till de mer genomgripande förändringar som har diskuterats .
då gives också tillfälle att finna nya gemensamma lösningar och analysera ändringsförslagen från utskottsdebatten .
rättstillämpningen i konkurrensfrågor måste vara korrekt .
felaktigt tillämpad konkurrenspolitik kan orsaka rättsförluster och göra ingrepp i äganderätten , vilket är en viktig , grundläggande princip som vi skall slå vakt om .
det ligger en ganska spännande debatt framför oss .
en konferens där frågorna ventileras möjliggör att missförstånd kan rätas ut , samtidigt som vissa punkter också kanske kan förbättras .
parlament och kommission kan tillsammans stärka insatserna för en effektiv konkurrenspolitik och därmed skapa nya möjligheter och nya resurser för medborgarna .
just i min valkrets , stockholm , har vi många goda lokala exempel på ökat utbud och förbättrad kvalitet som uppstått just på grund av konkurrensutsättningar på tidigare helt monopoliserade områden .
vi tillskyndar en fortsättning på den öppna debatt som stärkts under behandlingen av betänkandena av von wogau och rapkay .
vi hoppas att de rättsliga synpunkterna också kommer att tillmätas den vikt som är rimlig i en rättsstat .
herr talman , kära kolleger ! det gläder mig att jag får hålla mitt första tal här i dag som ny ledamot , även om det sker med en viss försening .
först vill jag tacka föredragandena von wogau , langen , rapkay , jonckheer samt kommissionen för det mycket goda samarbetet .
konkurrensen utgör säkerligen grundvalen för en marknadsekonomi med socialt ansvar , och den europeiska konkurrenspolitiken har varit framgångsrik , inte minst vad gäller energi och telekommunikation , och har lett till märkbart lägre priser och bättre service .
allt till konsumenternas fördel .
men nu har vi kommit fram till en punkt där vi måste vidareutveckla konkurrenspolitiken .
här har kommissionen lagt fram en ny vitbok med två kärnpunkter : anmälningsplikten skall överges , och den rättsliga verkställigheten skall återföras .
att man överger anmälningsplikten innebär i varje fall mindre byråkrati och administrativa kostnader .
denna systemändring leder naturligtvis samtidigt till mer ansvar för de enskilda i näringslivet .
det är inte längre så enkelt att man bara lägger fram något och får det godkänt , utan nu måste alla till att börja med själva bära ansvaret , och det är kanske också orsaken till att en eller annan där ute uppfattar detta som obehagligt .
men jag tror att vi bör utnyttja chansen att låta europa också ge en signal till mindre byråkrati .
den andra punkten är återföringen av den rättsliga verkställigheten .
för att en rättslig kultur skall kunna skapas i europa måste rätten givetvis inte bara tillämpas av kommissionen och av centrala organ , utan också av nationella myndigheter och domstolar .
vi säger ju inte heller att all eg-rätt alltid skall beslutas centralt , men just i anpassningsfasen kommer det att finnas en viss osäkerhet vad gäller rätten .
här är det säkerligen nödvändigt , i det lagstiftningsförfarande som vi står inför , att utveckla ett instrument för att ge företagen rättssäkerhet och möjlighet att vända sig till kommissionen .
det bör hållas en dörr öppen till en europeisk kartellmyndighet , som säkert kommer att diskuteras i framtiden .
men vi behöver mer öppenhet i konkurrenspolitiken .
parlamentet måste bli mer delaktigt , och jag tror också att om vi inför ett register , där vi kan se vilka statliga åtgärder som vidtas , så kommer detta att leda till disciplinering i medlemsstaterna .
vad gäller konkurrensen i framtiden ligger emellertid två punkter mig mycket varmt om hjärtat .
det ena är subsidiariteten .
vi anser alla att konkurrens är nödvändig för ekonomin och främjar prestationsförmågan , och jag tror att vi också bör släppa in konkurrens i regionerna .
konkurrensen mellan regionerna kommer säkerligen att stärka europeiska unionen , och inte försvaga den .
här kan jag nämna exemplen med ga-stöd , sparkassor och delstatsbanker , samt kvalitetsgaranti .
här har en region av egen kraft skapat något för att saluföra sina egna produkter .
dessa egna initiativ får inte förstöras från europeiskt håll .
jag tror att det också är nödvändigt med en höjning av deminimus-bestämmelserna .
vi bör satsa allt på att påskynda konkurrensen mellan regionerna .
det andra är en diskussion om konkurrens och marknadsekonomi med socialt ansvar , och då talar jag här inte om misslyckanden från marknadens sida .
jag har ju redan nämnt exemplen med delstatsbanker och sparkassor , men jag vill driva det som man alltid hör från det ena eller andra hållet till sin spets .
en boende på ett ålderdomshem är i dag socialt placerad .
men man kan också betrakta honom som en kund , och jag tror att vi ganska tydligt och i god tid bör diskutera var det sociala området , var de strukturer som vuxit upp sätter stopp för konkurrensen .
annars kan jag här använda uttrycket kunder för detta område , och därigenom mycket starkt förstöra sociala områden .
slutligen vill jag också säga i fråga om subsidiaritetsprincipen : jag anser att det är absolut nödvändigt att där medlemsländerna medger att regioner och kommuner kan uppbära skatter skall detta bibehållas och inte regleras enhetligt av europa .
. tack så mycket , herr kollega .
jag gratulerar er till det som man inom den tyska parlamentarismen , i ert fall felaktigt , kallar för ett jungfrutal .
herr talman , herr kommissionär , kära kolleger ! jag kommer att tala å min kollega robert goebbels vägnar , eftersom han inte kunde komma på grund av politiska förpliktelser .
inom utskottet för ekonomi och valutafrågor väckte jonckheerbetänkandet bittra kontroverser kring marknadens sätt att fungera .
en knapp högermajoritet lyckades stryka samtliga hänvisningar till att marknaden har brister .
men även om majoriteten i vårt parlament skulle följa denna ultraliberala uppfattning om en så kallad perfekt marknad , skulle världen inte förändras för det .
ekonomiska rapporter från den verkliga världen ger tillräckliga bevis för att man inte på något sätt skapar en perfekt konkurrens och bästa möjliga resursfördelning genom att avskaffa alla former av offentliga interventioner på marknaden .
marknaden må ha varit människors främsta handelsplats sedan urminnes tider , men den har aldrig varit perfekt .
marknaden gynnar kortsiktighet och omedelbara vinster .
på marknaden verkar styrkeförhållandena mellan utbud och efterfrågan i allmänhet till de svagares nackdel , konsumenterna , arbetarna .
för att fungera fordrar marknaden regler .
den nödvändiga och värdefulla initiativandan måste åtföljas av en känsla av ansvar gentemot samhället .
vi europeiska socialister är för en marknadsekonomi med sociala ändamål .
marknaden är inte ett mål i sig ; den skall bidra till att förbättra de mänskliga villkoren .
europeiska unionen och staterna skall inte ta de ekonomiska aktörernas plats , men statsmakterna måste fastställa regler och mål som gör att ekonomin kan utvecklas på ett hållbart sätt .
statliga stöd kan slutligen möjliggöra omstruktureringar , erbjuda utbildning , rädda arbetstillfällen och därmed kunnande .
huvudmålet med unionens konkurrenspolitik får inte vara att minska den allmänna stödnivån .
de statliga stöden måste anpassas efter unionens mål , framför allt ekonomisk och social sammanhållning , hållbar utveckling samt forskning .
kommissionen måste bedriva klappjakt på illegala stöd och de stöd som verkligen blockerar den inre marknaden .
men att avskaffa alla former av statsstöd skulle vara ett allvarligt misstag .
internet är inte en marknadsprodukt , utan resultatet av forskning som finansierats av den amerikanska armén .
world wide web , som har möjliggjort en blixtrande utveckling av informationssamhället , utvecklades av europeiska atomforskningscentret ( cern ) i genève , återigen med hjälp av statsstöd .
att den tyska regeringen räddade holzmann-gruppen kritiserades som ett ogrundat hinder mot marknadsekonomin .
centralbankschefen duisenberg försökte till och med skylla eurons svaghet gentemot dollarn - för övrigt tämligen relativ - på denna statliga interventionism .
jag har inte hört duisenberg kritisera det faktum att de amerikanska penningpolitiska myndigheterna räddade hedge fund ltcm .
att vilja rädda 60 000 arbetstillfällen , det är uppenbarligen att begå en synd gentemot marknaden , men att rädda kapital tycks inte skapa några problem för den fria marknadens förespråkare .
man uppbringar offentliga medel för att reparera de skador som har orsakats av den internationella spekulationen , bl.a. i mexiko , asien och brasilien .
människors arbete betraktas däremot som vilken justeringsfaktor som helst .
vi socialister avvisar denna liberala världsfrånvända inställning .
vi vill ha en riktig konkurrenskultur i europa .
den statliga handen måste förbli synlig för att styra marknaden , och kommissionen bör vara dess domare .
herr talman , bästa kommissionär och kära kolleger ! jag vill börja med att tacka herr rapkay för ett väl utarbetat betänkande och ett gott samarbete .
kommissionär monti ! jag vill tacka er för ett utmärkt samarbete och jag vill säga till er att ni nu vid årtusendeskiftet har en mycket viktig funktion .
ni skall ju städa upp efter de nationella regeringar som har stora visioner på konkurrenspolitikens område , men endast fantasin sätter gränser för vilka olyckor de nationella regeringarna kan åstadkomma .
jag kan här nämna de senaste exemplen vi har sett : holzmann , ett företag som fått ett omfattande stöd från den tyska regeringen , sågverk i f.d. östtyskland och inte minst stöden till skeppsvarven .
detta är tre områden inom vilka många danska företag har stora problem och blir utkonkurrerade från marknaden .
jag vill säga till herr poos att jag är helt överens med ordförande duisenberg om att det finns exempel på att några av europeiska unionens medlemsstater inte är förmögna att omstrukturera sina ekonomier , och därmed bidrar till att undergräva eurons värde .
den liberala gruppen har lagt fram 80 ändringsförslag i utskottet , som alla rör statligt stöd .
det är förslag som vi anser leder fram till genomblickbarhet och öppenhet , vilket är mycket viktigt när det gäller att få den inre marknaden att fungera .
jag vill gärna ta tillfället i akt och tacka mina kolleger i utskottet för deras stöd till den liberala gruppens förslag .
våra förslag rör som sagt möjligheten till insyn , och jag vill gärna betona det ändringsförslag som uppmanar kommissionen till att utarbeta enhetliga kriterier och villkor för den typ av statligt stöd som vi anser vara lagligt , just för att se till så att företagen kan planera sin situation .
en annan sak är frågan om vad vi skall göra om det statliga stödet förklaras olagligt .
hur ser vi till att få det olagligt utbetalade statliga stödet tillbaka ?
i dag finns inga gemensamma bestämmelser på detta område och vi uppmanar kraftfullt kommissionen att skapa en harmonisering av bestämmelserna om återbetalning .
detta är enda sättet för att säkerställa enhetliga konkurrensvillkor .
till sist föreslår vi att vi dels skapar ett register , vilket flera av mina kolleger varit inne på , men också en resultattavla som visar var länderna står i dag vad gäller statligt stöd .
ni har visat oss vägen , herr monti , med en resultattavla för den inre marknaden .
det är detta som inspirerat oss till att föreslå samma sak vad gäller statligt stöd .
jag hoppas verkligen att kommissionär monti kommer att stödja dessa förslag , och jag ser fram emot era kommentarer och er ståndpunkt .
avslutningsvis vill jag hälsa kommissionens xxviii : e rapport om konkurrenspolitiken välkommen ; ännu en gång får vi ta del av ett väl utfört arbete .
men som jag redan har nämnt bör det övergripande syftet fortfarande vara genomblickbarhet och öppenhet .
det finns fortfarande behov av en uppryckning inom de nämnda områdena och det finns därför en god anledning till att fortsätta med att arbeta på ett målinriktat sätt för att lösa problemen rörande den bristande genomblickbarheten och öppenheten på området för statligt stöd .
det är inte minst nödvändigt i förhållande till den kommande utvidgningen , och jag vill gärna tacka herr jonckheer som i sitt betänkande mycket grundligt behandlar problemen i samband med utvidgningen och hur vi skall se till att dessa länder uppfyller våra krav , men också hur vi säkerställer lika konkurrensvillkor .
det är klar att vi som liberala och gröna har olika uppfattningar om hur vi vill att världen skall se ut , men vad gäller vår målsättning är vi i stort sett överens , och vi vill försöka hitta en förnuftig lösning på våra problem .
herr talman , herr kommissionär ! vi har egentligen endast två frågor att svara på .
är statliga företagsstöd och avtal mellan företag legitima i en marknadsekonomi ? och : vem skall kontrollera undantagen till marknadsekonomins absoluta regler ?
på den första punkten vill vi mycket klart och tydligt säga att det i vissa fall krävs statliga företagsstöd , om vi skall ta hänsyn till de krav på en hållbar utveckling som europeiska unionen skriver under på , och det oavsett om det sker i form av skattelättnader , differentierad beskattning eller helt enkelt direkta stöd .
det är också berättigat att det skall kunna finnas avtal och begränsningsavtal mellan företag , eftersom alla sådana avtal bidrar till att dämpa konkurrensens negativa bieffekter på det sociala och miljömässiga planet .
vi svarar alltså mycket klart och tydligt ja - statliga stöd och avtal är legitima , men vi menar också att varje avtal verkligen måste åtföljas av en motivering .
i von wogaubetänkandet föreslår man att kontrollen av legitimiteten skall återföras till nationell nivå .
för oss förefaller det ganska riskfyllt , men vi kommer ändå att rösta för , eftersom vi medger att kommissionen inte kan göra allt .
vi kräver största möjliga öppenhet och att kommissionen skall anförtros största möjliga undersökningsmakt för att i efterhand kontrollera om beviljade undantag är legitima .
herr talman ! ännu en gång diskuterar vi europeiska unionens konkurrenspolitik .
men under vilka förhållanden förs denna debatt , och vilka slutsatser bör vi komma fram till ?
dagens verklighet kännetecknas av gigantiska fusioner och sammanslagningar av enorma monopolföretag och skapandet av världsomspännande koncerner med fruktansvärd makt .
borde vi inte ta upp detta i vår debatt ?
vilken konkurrenspolitik vill och kan införa kontroller av dessa monopolföretags verksamhet ?
vissa branscher inom den europeiska industrin , t.ex. varvsindustrin , flygtransporterna , stålindustrin , har drabbats enormt hårt av den konkurrenspolitik som bedrivs .
de har förlorat viktiga marknadsandelar inom världshandeln och hundratusentals arbetstillfällen .
skall vi inte ta upp detta till diskussion ?
den skandalösa maktkoncentrationen inom strategiskt viktiga sektorer gör att vinstinriktade multinationella företagsgrupper får kontroll över ekonomin i hela länder - även i unionens medlemsländer .
trots detta envisas vi med en fortsatt försvagning av den offentliga sektorn , och vi är beredda att skärpa konkurrenspolitiken ytterligare , när vi anser att statliga beställningar från företag av offentlig karaktär också är ett slags statligt stöd .
å andra sidan leder bortfallet av hundratusentals arbetstillfällen till en våldsam ökning av arbetslösheten .
arbetstagarna utsätts för ett enormt angrepp på sina arbetsrättsliga och sociala rättigheter .
konsumenterna ser hur deras levnadsstandard sjunker , hur fattigdomen breder ut sig och hur den offentliga sektorn och den produktiva basen i de flesta av unionens länder skärs ned och upplöses till förmån för en ohämmad och fördärvbringande konkurrens , den totala marknadsekonomin och storkapitalets monopolintressen .
jag anser att det även är den förda konkurrenspolitiken som bär ansvaret för allt detta , och jag tar fullständigt avstånd från den .
herr talman , herr kommissionär ! under brytningsåret , före övergången till den gemensamma valutan , gjorde kommissionen stora ansträngningar för att euron skulle kunna införas under gynnsamma omständigheter .
konkurrenspolitiken bidrog till denna tilldragelse , inom ramen för dessa medel .
vi är för vår del fortfarande bestämda motståndare till den gemensamma valutan , som långt ifrån ger oss fördelarna och flexibiliteten med en gemensam valuta , utan i stället stänger in oss i en artificiell tvångsstruktur som påtvingats europas folk .
men att styra är samtidigt att förutse och även att ta ansvar , och i det nya framtvingade sammanhanget spelar konkurrensrätten naturligtvis en viktig roll .
på det området har kommissionen prioriterat flera handlingslinjer : att påverka marknadernas struktur genom att aktivt motverka konkurrenshämmande metoder , att inrikta kontrollverksamheten på de affärer som har ett uppenbart gemenskapsintresse samt att markera sin önskan om en modernisering av konkurrensrätten .
vad gäller statliga stöd måste man se till att bestämmelserna inte blir för tungrodda . enligt vår uppfattning är det därför inte önskvärt att införa ett offentligt register över samtliga stöd , eftersom denna tyngande förpliktelse givetvis skulle gå på tvärs mot försöken att lätta på de byråkratiska kraven .
när det slutligen gäller en modernisering av tillämpningen av artiklarna 85 och 86 i fördraget , anser vi inte att en decentraliserad tillämpning nödvändigtvis är ett steg i rätt riktning .
kommissionen skulle inte endast behålla sin makt att undanhålla de nationella myndigheterna ett ärende - de nationella domstolarna har också klara förpliktelser att undvika varje form av konflikt med kommissionens beslut .
nationalstaterna skulle således bli kommissionens världsliga rättvisa , med uppdraget att garantera en respekt för tillämpningen av regler som de inte har någon kontroll över .
sammanfattningsvis vill jag säga att även om vissa bestämmelser går i rätt riktning , kommer vi självklart att förbli vaksamma för att förhindra en federalistisk utveckling , vilket skulle skada europa och staternas suveränitet .
herr talman , herr kommissionär , ärade kolleger ! vi är i allt väsentligt positiva till kommissionens vitbok om konkurrensen , framför allt när det gäller avskaffandet av systemet med meddelande och tillstånd , men vi är också en aning frågande inför ett par punkter .
framför allt finns risken att delegering av behörigheter till de enskilda staterna , något som i flera avseenden är nödvändigt , kan leda till en alltför kraftig expansion av konkurrensinitiativen och att någon kan frestas att använda antitrustbestämmelserna , inte som en yttersta garanti för att marknaderna skall fungera väl och så som var avsett , utan som ett instrument för den egna ekonomiska och industriella politiken , som ett instrument för planering och ingrepp i marknadernas egna spontana dynamik eller kanske till och med som ett verktyg för protektionistisk politik .
i det avseendet tror jag att vi kan finna vägledning i det som von eieck har skrivit och säkerligen också i det som den store italienske liberalen bruno leoni säger när han just varnar för riskerna för en kraftig ökning av konkurrenshämmande åtgärder .
det allvarligaste hotet mot marknaden , konkurrensen och valfriheten för de europeiska användarna och konsumenterna är fortfarande hotet om statliga ingrepp i ekonomin .
det finns statliga stöd till företagen , det har vi redan talat om , det finns fortfarande en stark offentlig närvaro i ekonomin - tänk till exempel på att det italienska finansdepartementet kontrollerar 15 procent av allt kapital på italienska börsen - det finns hinder som regeringar och centralbanker reser inför verksamhet som innebär merger and acquisition ; vi har ofta under de senaste dagarna hört talas om fallet vodafone-mannesmann och räddningen av osman .
slutligen , herr kommissionär , får vi inte glömma att det fortfarande finns stora ekonomiska sektorer som är i offentliga händer , från den statliga televisionen , som tvångsfinansieras av licensinnehavarna , och postverken , till vissa obligatoriska försäkringssystem , inklusive sjukvårds- och olycksfallsförsäkringar , som hanteras av ineffektiva offentliga monopol som inte ger något val åt användarna om de inte är mycket välbeställda .
herr kommissionär , jag känner väl till fördragets begränsningar , men jag anser att det även i detta fall är viktigt att understryka att den europeiska ekonomin drabbas hårt av konkurrensen från den amerikanska , även och framför allt på grund av bristen på möjligheter och konkurrens .
det som vi gör här är förmodligen mycket viktigt , men det är fortfarande otillräckligt .
herr talman ! vi för en speciell debatt : om konkurrenspolitik och om statsstöd , statens vänstra och högra hand så att säga .
medan emu-kriterierna tvingar medlemsstaterna att begränsa sina utgifter har den höga nivån i fråga om statligt stöd till företagslivet kvarstått .
förståeligt , för den medlemsstat som börjar med att avveckla statligt stöd löper den största risken att drabbas av företag som flyttar ut , med negativa följder för sysselsättningen .
men samtidigt obegripligt , för dålig företagaranda och icke livsdugliga arbetsplatser skall inte understödjas med pengar från skattebetalarna .
i princip är enbart horisontala åtgärder tillåtliga eftersom de inte eller knappast rubbar konkurrensen .
föredragandens ändringsförslag 6 och 7 förtjänar därför stöd .
ändringsförslagen 1 och 5 visar på fenomenet att marknaden inte fungerar , för enbart marknadsinstrumentet leder inte till det ideala samhället .
det är de sårbara människorna som befinner sig i det hörn där motgångarna slår .
marknadsverkan måste användas på ett listigt sätt för att låta medborgarnas och företagens ansvar komma till sin rätt maximalt .
om denna ansträngning misslyckas måste en statsmakt ingripa .
kommissionens vitbok om modernisering av konkurrenspolitiken liknar mer ett diskussionsdokument .
pläderingen för decentralisering för att lätta arbetsbördan inom generaldirektoratet för konkurrens ger ett sympatiskt intryck , men det sätt på vilket kommissionen vill utforma denna tanke leder till att den rättsliga makten blir överbelastad .
det går ut över rättssäkerheten för näringslivet .
minskar verkligen kommissionens arbetsbörda när nationella domstolar är skyldiga att rapportera till kommissionen ?
vilken åsikt har rådet om detta , och är kommissionären beredd till en grundlig omprövning av dessa punkter ?
en vitbok är definitionsmässigt inte något som man tar till sig eller lämnar därhän ; den syftar till att väcka reaktioner , och det har denna vitbok helt klart lyckats med .
den utgör ett gott diskussionsunderlag , och i den bemärkelsen är den välkommen .
jag förstår författarnas utgångspunkter och stöder dem .
jag utgår också från att ni , herr kommissionär , vill värna om era företrädares rykte och det de byggt upp , och att era tjänstemän har samma mål .
jag kan inte föreställa mig att kommissionen skulle ta initiativ till att inleda en grundlig aveuropeisering eller till att börja åternationalisera . men jag känner ändå en viss oro , ändå har jag frågor .
för det första gäller det sammanhållningen då politiken skall omsättas i praktiken .
allmänt sett är jag en stark förespråkare för kulturell mångfald , men inte på området konkurrenskultur på den inre marknaden .
den inre marknaden behöver en enhetlig konkurrenspolitik , inte bara vad konceptet beträffar , utan även i fråga om att omsätta den i praktiken .
det kommer visserligen europeiska förordningar och tolkningsmeddelanden .
kommissionen borde också ha rätt att ta upp ärenden och ge riktlinjer åt de nationella konkurrensmyndigheterna .
men jag ställer mig ändå frågan om vi inte löper risken att hamna i en långdragen process , där vi hela tiden skulle bli tvungna att ta ett steg tillbaka innan vi kan ta två steg framåt .
jag skulle således vilja veta mer , herr kommissionär , om på vilket sätt kommissionen kommer att garantera en enhetlig omsättning i praktiken och om ni själv anser att de vägar som skisseras från och med punkt hundra i vitboken är genomförbara .
för det andra förstår jag näringslivets oro i fråga om rättssäkerheten .
nu anmäls många ärenden just med tanke på detta .
i framtiden bortfaller detta instrument .
i vitboken säger ni att kommissionen ändå kommer att fatta individuella beslut som kan tjäna som riktlinjer , men vilka kriterier kommer ni att tillämpa för att den ena gången fatta ett sådant beslut och den andra gången inte ?
för det tredje vill jag gärna veta om kommissionen har undersökt vilka konsekvenser dess nya tillvägagångssätt kommer att få för näringslivets strategi .
jag är särskilt oroad över de små och medelstora företagens öde , vilka förlorar ett visst juridiskt och ekonomiskt skydd i likhet med vad som måste vara fallet i fråga om det nya gruppundantaget för distributionssektorn .
för det fjärde skulle jag gärna vilja veta varför kommissionen inte beslutat sig för att låta nullitetssanktionen träda i kraft ex tunc då det rör sig om tydliga överträdelser av konkurrensreglerna .
för det femte handlar det om den utvidgning som står för dörren , och jag frågar mig om kandidatländerna kommer att kunna mäkta med att spela vårt spel .
i själva verket ligger de fortfarande i träning .
vilka garantier har vi för att de kommer att växa ut till förstaklasspelare i den interna marknadens liga ?
för det sjätte och sista påminner jag om en punkt som jag också tog upp i mitt betänkande om de vertikala restriktionerna , i synnerhet företagsjuristernas så kallade legal privilege .
om kommissionen genomför sina föresatser i vitboken förefaller det mig som om diskrimineringen på den inre marknaden mellan de externa och de interna juridiska rådgivarna kommer att bli större och således också mer oacceptabla .
överväger kommissionen att göra något för att bevilja företagsinterna jurister i alla medlemsstater ett legal privilege ?
herr kommissionär ! jag ställer dessa frågor som försvarare av den inre marknaden , och jag hoppas att vi här i den bemärkelsen allesammans är partner och att diskussionen mellan dessa partner inte kommer att bli steril utan kommer att kunna bära frukt .
herr talman ! jag vill inleda mitt anförande om vitboken med att framföra mina gratulationer till föredragande von wogau .
ett tydligt bevis på den höga grad av enighet som råder mellan europeiska socialdemokratiska partiets grupp och hans betänkande är att endast ett ändringsförslag har lagts fram under ärendets gång .
vi ställer oss således positiva till betänkandet , precis som vi ställer oss positiva till de grundläggande inslagen i vitboken , herr kommissionär .
gemenskapens konkurrensbestämmelser har , ända sedan fördraget trädde i kraft , varit en av gemenskapspolitikens grundvalar .
efter nästan fyrtio år i kraft har dessa bestämmelser börjat visa sig vara föråldrade .
därför är det angeläget med en modernisering .
denna modernisering är nödvändig i synnerhet på fem punkter .
punkt ett : systemet för godkännande ; punkt två : den decentraliserade tillämpningen ; punkt tre : bestämmelserna för förfarandena ; punkt fyra : rättstillämpningen och slutligen punkt fem : paragrafrytteriet .
det har funnits ett överhängande behov av en reform av systemet för enstaka beviljanden , och en sådan har enhälligt efterfrågats av företag , forskare och advokater med specialistkompetens .
jag har inte deltagit i en enda sammankomst för experter på gemenskapens konkurrensbestämmelser , där man inte har begärt en ändring av systemet .
ett system som medger så pass få beslut , i form av beviljanden eller förbud , som det nu rådande systemet är inte godtagbart .
artiklarna 81.1 och 82 har sedan länge kunnat tillämpas av de nationella konkurrensmyndigheterna .
däremot har man inte kunnat tillämpa artikel 81.3 , något som i viss mån har förhindrat en följdriktig tillämpning av artikel 81.1 .
för närvarande har , som mina damer och herrar vet , två tyska domstolar vardera anhängiggjort ett mål för förhandsavgörande vid eg-domstolen , med ifrågasättanden av om det är möjligt att tillämpa artikel 81.1 då artikel 81.3 inte kan tillämpas .
därför är en reform på den punkten oumbärlig .
grunderna för konkurrensförfarandet fastslås i förordning nr 1762 .
man röstade enhälligt för en ändring .
det faktum att förordningen inte fastslår ett regelrätt förfarande , inte fastställer några tidsramar , inte reglerar de inblandade parternas tillgång till handlingarna och inte på ett relevant sätt erkänner rätten till försvar , har varit motiv till det enhälliga kravet på en reform .
eg-domstolen har för länge sedan godtagit att gemenskapens konkurrensbestämmelser tillämpas av medlemsstaternas rättsskipande organ , och kommissionen offentliggjorde redan 1994 ett meddelande i den frågan .
således är det nödvändigt att underlätta ett sådant förfarande .
paragrafrytteriet är något av det som starkast kritiseras i gemenskapens konkurrensbestämmelser .
bedömningen av om vissa avtal är konkurrensbegränsande eller ej beror , till följd av den kontinentala rättstraditionen , snarare på en analys av avtalets klausuler än av effekten på marknaden .
av den anledningen har det varit nödvändigt att inbegripa en ekonomisk analys .
genom vitboken försöker man lösa dessa problem , och därför stöder vi förslagen i denna .
vi har även upptäckt vissa brister i betänkandet .
bland dessa kan i första hand nämnas att man , trots att det handlar om en modernisering av artiklarna 81 och 82 , lägger hela tyngdpunkten på artikel 81 och inte på artikel 82 .
i en tid då processer med samordning av företag , eller privatiseringen av monopol intar en framskjuten och till med förstärkt ställning , är det särskilt viktigt att motarbeta orimliga förfaranden .
för det andra bör förordning nr 1762 upphävas och ersättas med en ny förordning .
på den punkten stöder vi betänkandet .
skulle däremot några av ändringsförslagen godkännas , och då i synnerhet de som framlagts av europeiska folkpartiets grupp , anser vi att betänkandet förvanskas , att det förvandlas till ett motsägelsefullt dokument utan stringens , och i sådant fall kommer vi att bli tvungna att ompröva vårt stöd .
herr talman , mina damer och herrar ! bland alla de frågor som diskuteras i denna gemensamma debatt , vill jag koncentrera mig på några tankar kring det vår kollega berenguer talade om , det vill säga den modernisering av konkurrenspolitiken som åsyftas i kommissionens vitbok .
jag anser uppriktigt sagt att denna modernisering är tillfredsställande .
kommissionär monti har uppnått goda resultat i sitt arbete , precis som sin föregångare , och har tydligt visat att han , vid sidan av skapandet och utvecklandet av en inre europeisk marknad , haft förmåga att vidta de rätta åtgärderna för att marknadsekonomin inom unionen skall fungera , utan de avvikelser som vi ekonomer vet kan förekomma i samband med att marknaden expanderar , på det sätt som den har gjort inom europeiska unionen sedan 1993 .
om allting fungerar , om vi är nöjda , om kommissionens agerande i huvudsak har varit korrekt , varför behövs det då en ändring ?
olika argument har lagts fram som talar för detta .
berenguer har gjort en högst korrekt analys , där han visar på behoven och reformerna till följd av dessa i syfte att förbättra konkurrenskraften , men jag finner det angeläget att man garanterar att den standard och de kriterier som tillämpas av respektive myndighet i medlemsstaterna överensstämmer i alla avseenden .
för om de inte gör det , hamnar vi i en paradoxal situation , där kommissionen själv är den som inför illojala konkurrensmedel på den inre europeiska marknaden .
i sådana fall har vi inte gjort några framsteg , utan det skulle tvärtom innebära att vi gick bakåt i vår tillämpning av konkurrenspolitiken inom unionen .
herr talman ! till att börja med vill jag uttala mitt erkännande till kommissionen för den förbättring som den xxvii : e rapporten om konkurrenspolitiken i unionen innebär i förhållande till tidigare utgåvor .
likaså vill jag framhålla det arbete som har utförts av föredragande rapkay , som har gjort en kort och koncis analys av en så pass tjock och omfattande text som denna .
jag stöder helt hans påpekande om behovet av att ge handlingsutrymme åt regioner - som till exempel baskien som jag själv företräder - till följd av subsidiaritetsprincipen .
ändå kan jag inte glömma den kritik som vid flera tillfällen har framförts , såväl av medlemsstaterna som av marknadsaktörerna som , utifrån det begränsade handlingsutrymme , den begränsade valfriheten som kommissionen har när den skall bedöma varje enskilt fall , hävdar att det rättsliga läget är osäkert , eftersom det inte finns några tydliga spelregler som gör att de inblandade kan förutse myndighetens ställningstagande och utifrån det göra korrekta ansökningar om bidrag till främjande åtgärder för den ekonomiska verksamheten och sysselsättningen , förslag om sammanslagning av bolag , etc.
det enda säkra sättet har blivit att begära ett godkännande i förväg , via enskilda ärenden där det dröjer minst sex till åtta månader innan besked lämnas , en alldeles för lång tidsperiod som endast åtföljer problemen med bristande rörlighet till sådan verksamhet som genererar välstånd och sysselsättning .
jag tycker att det saknas , och föreslår av den anledningen , att man fastställer ett flertal bestämmelser , tillkännager tydliga spelregler som vi alla har att vinna på : företagare , investerare , arbetstagare och befolkningen i allmänhet .
herr talman , parlamentskolleger ! jag vill gärna understryka att i en period av stora tekniska förändringar - se bara på det som sker inom informationstekniken eller inom andra sektorer som energi och transporter - är skyddet av konkurrensen av grundläggande betydelse för vår framtid .
när det gäller den ekonomiska tillväxten , och därmed ökningen av sysselsättning och välfärd , blir skyddet av en konkurrensfrämjande politik i våra länder inom unionen en avgörande faktor av grundläggande betydelse för vår framtid .
det är av den anledningen jag uttrycker mitt starka stöd för den här aktuella betänkandet .
jag har noterat att kommissionen under den senaste perioden har ansträngt sig för att hävda den principen kraftfullt och entydigt , just för att skydda marknadernas flexibilitet , såväl marknaderna för produkter som för tjänster .
jag hävdar bestämt att detta kommer att vara av yttersta vikt för vår framtid , för den europeiska ekonomin och framför allt för att skydda vårt välstånd och den allmänna tekniska utvecklingen i europa .
herr talman ! för de konservativa i storbritannien är tillämpningen av den europeiska konkurrenspolitiken på ett effektivt och enhetligt sätt kärnfrågan när det gäller att skapa en effektiv inre marknad i hela europeiska unionen .
därav följer att alla förslag som innebär större förändringar av systemet för att genomdriva konkurrenspolitiken måste granskas ingående och noggrant .
sanningen är att den inre marknaden ännu inte är fullständig .
under mina sex månader som ledamot av detta parlament har jag blivit mycket medveten om många ledamöters beslutsamhet att driva det som beskrivs som det europeiska projektet framåt .
dagligen hör vi talas om behovet att verka för ett vidare och djupare europa .
men allt detta är i realiteten bara retorik när vi tittar på de nationella , regionala och lokala hinder som fortfarande står i vägen för en sann europeisk inre marknad .
det är i detta sammanhang jag vill se kommissionens förslag .
jag skulle vilja göra klart att vi har det största förtroende och respekt för kommissionär monti .
vi ser honom som mannen som skall utrota karteller .
men han skulle förstå att vi , liksom med alla andra , måste bedöma hans enskilda förslag och underkasta dem en grundlig granskning .
detta är vad vår föredragande i utskottet för rättsliga frågor och den inre marknaden , von wogau , har gjort .
jag vill gratulera honom , tråkigt nog i hans frånvaro , till det grundliga och noggranna sätt på vilket han har sammanställt detta betänkande - och också för att han har stått ut med att jag har varit så besvärlig !
han nämnde tidigare att betänkandet antogs med en betydande majoritet , men inte med mitt stöd .
så även om jag inte delar hans slutsatser anser jag att han i sitt betänkande har belyst många av de frågor kommissionen måste ta upp .
den första är möjligheten att åter göra konkurrenspolitiken till en nationell fråga .
jag vet att kommissionen är negativ till detta , men möjligheten finns .
jag är fortfarande orolig över nationella domstolars och konkurrensmyndigheters kapacitet .
jag är fortfarande orolig över hur den rättsliga processen som helhet fungerar .
härom dagen frågade jag kommissionär monti vad som händer om han har fel och konkurrenspolitiken i praktiken åter blir nationell .
von wogau sa att vi kan titta på eg-domstolen .
vi i storbritannien tittar just på eg-domstolen för tillfället .
vi finner då att eg-domstolen inte klarar av att ge oss interimsåtgärder för en viss tvist vi har med frankrike för ögonblicket , och där vi har kommissionens stöd .
för att ingen skall tro att detta bara är en nationell fråga tog det tio år för eg-domstolen att döma i factortame-fallet , där den brittiska regeringen var den svarande .
så någonting måste göras åt rättsskipningen .
jag frågar kommissionen vad som kan göras för att snabba upp tillämpningen på detta speciella område .
vad gäller visshet om rättsläget instämmer jag i thyssens poäng .
det är viktigt att företagen har visshet om rättsläget .
jag nämnde detta för kommissionär monti igen nyligen .
han sade att vi inte alltid får låta oss ledas av advokater .
jag måste säga att jag berörs av detta som advokat men också som tidigare konkurrensminister i storbritannien .
vi har ju alla vårt förflutna att dras med , men det är viktigt att företagen har visshet om rättsläget .
jag skulle också vilja fråga kommissionen om den har analyserat hur denna förändring påverkar industrin : en samhällsekonomisk kostnads-intäktsanalys av det slag som nu håller på att bli en del av den europeiska politiken .
jag vet att det har gjorts en analys av hur kommissionen påverkas av förändringen .
vi har fått veta att människors tid slösas bort för närvarande och att förändringarna därför skulle kunna vara till fördel .
men jag anser verkligen att vi under dessa omständigheter behöver veta vilken inverkan de får på företagen .
slutligen söker vi som brittiska konservativa en ändrad inriktning , mot skapandet av en oberoende konkurrensmyndighet .
jag skulle vilja höra vad kommissionär monti har att säga om det .
herr talman ! alltsedan den europeiska integrationen började har europeiska unionens konkurrenspolitik varit av central betydelse .
den kan indelas i spänningsförhållandet , som också innefattar konceptet för den europeiska integrationen , solidariteten mellan medlemsstaterna , samarbetet mellan medlemsstaterna för att utforma bättre och mer effektiva ramvillkor för människorna och näringslivet , och konkurrensen som skall skapa impulser för att förbättra europeiska unionens konkurrenskraft och förmåga inför framtiden .
konkurrenspolitiken är därför med all rätt ett av de viktigaste politiska områdena .
vi kan vara stolta över att ha en europeisk konkurrenskultur som också faktiskt syftar till att genomföra en marknadsekonomi med socialt ansvar .
vi kan vara stolta över kartell- och fusionskontrollen .
men vi måste vara vaksamma när det gäller de aktörer som verkar över hela världen , som det nationella agerandet inte längre kan sätta några gränser för .
man måste tänka på en ordvändning hos den franska författaren vivienne forestier , som beskriver tillståndet i världen som en ekonomins terror .
samhället överlämnar sig åt marknaden .
så vill vi inte ha det i europeiska unionen .
i en tidsålder av strategier rörande allianser och millenniefusioner - 1998 utbetalades 2 400 miljarder usd för övertaganden - vet vi att en konkurrensskadlig praxis stävjas inte bara med hjälp av våra egna bestämmelser , utan också via bilateralt samarbete med usa eller japan eller andra , så länge det fortfarande inte finns någon internationell konkurrensrätt , som absolut borde finnas !
europeisk konkurrenspolitik - detta glömmer vi ofta bort - är inte bara av betydelse för den rättvisa konkurrensen som sådan , utan också för prisutvecklingen , tillväxten och sysselsättningen och därmed också för medborgarna .
liksom de andra kollegerna kräver jag medbeslutande från europaparlamentet när det gäller konkurrensrätten .
det måste äntligen genomföras !
det är också viktigt att framhäva sammanhanget mellan konkurrenspolitik och konsumentskydd .
det är positivt att kommissionär monti på detta område vill uppnå framsteg i dialogen med europaparlamentet , men också i dialogen med de icke-statliga organisationerna , konsumentskyddsorganisationerna och medborgarna .
större öppenhet kommer också att bidra till en offentlig acceptans av konkurrenspolitiska beslut .
då kan man nämligen förstå , att exempelvis de lägre el- och telekommunikationspriserna också är ett resultat av den europeiska konkurrenspolitiken och att bryssel inte bara måste ställas vid skampålen när det fattas beslut om stöd , som i en aktuell eller lokal situation säkert kan förorsaka problem .
det måste också finnas klarhet särskilt om konkurrensreglerna med tanke på utvidgningen av eu .
det måste då framhävas att en statlig stödpolitik - detta framgår också tydligt av jonckheers betänkande - även i fortsättningen måste ge varje stat friheten att självständigt definiera och utforma sina offentliga uppgifter och ägandeförhållanden .
det måste därvid stå klart att stöden kan ha en nyttig funktion för att utjämna misslyckanden på marknaden och främja gemenskapens mål .
ett påpekande om vitboken : revideringen av artiklarna 81 och 82 innebär en vändpunkt i fråga om kartellbestämmelserna .
jag vänder mig mot detta , i motsats till majoriteten i denna kammare och även till majoriteten i min egen grupp , eftersom jag anser att systemet med direkt tillämplighet av undantagsregeln konkurrenspolitiskt är klart underlägset ett system där man har förbud med administrativt förbehåll , och därför att jag ser risken för en åternationalisering .
det rådande systemet medger öppenhet och erbjuder rättssäkerhet för företagen ; dess anmälningsplikt har utan tvivel lett till disciplinering och avskräckning .
problemet med för stor arbetsbörda som av kommissionen ställs i förgrunden är inte någon tillräcklig anledning till en djupgående ändring av rättssystemet .
här måste man också fråga sig om det över huvud taget kan genomföras utan en ändring i fördraget .
herr talman ! jag är mycket glad att randzio-plath nämnde den mycket viktiga bakgrunden till vår debatt , eftersom ingen talare hittills har gjort det .
eurons tillkomst i början av förra året släppte lös en enorm konkurrenskraft inom den europeiska industrin vilken bemöts av en sammanslagningsvåg av aldrig tidigare skådade proportioner .
till exempel visar nu siffrorna för förra året att det totala värdet av fusioner inom europa var 1,4 triljoner euro , vilket är sju gånger så mycket som vid höjdpunkten för den senaste europeiska fusionshaussen 1990 .
detta ställer konkurrenspolitiken inför enorma utmaningar , vilka jag hoppas att den kommer att leva upp till , eftersom många av dessa sammanslagningar helt visst kommer att vara utformade för att skydda företagens vinstmarginaler mot konkurrens snarare än att enbart stärka produktiviteten och ge dessa företag förmåga att verka i större skala .
kommissionär monti och hans kolleger står inför en ofantlig utmaning och eldr-gruppen är angelägen om att konkurrenspolitikens framstötar inte försvagas vare sig vad gäller granskningen av fusioner eller övervakningen av kartell- och monopolfrågor .
visst kan man delegera till nationella myndigheter , men vi skulle då vilja betona vad von wogau sade i sitt betänkande om behovet av en regelbunden övervakning av de nationella myndigheterna för att se till att det europeiska maskineriet inte slirar och speciellt be kommissionären att försäkra oss om att det dessutom kommer att förekomma stickprovskontroller .
herr talman ! jag vill under den korta talartid som står till mitt förfogande uttala mitt stöd för det arbete som har lagts ned av samtliga föredragande och även stödja mycket av det som här har sagts , i synnerhet av min kollega jonckheer , som kritiserar den alltför omfattande sammanställningen av fakta och påpekar behovet av insyn och av en socioekonomisk balans vad stödet beträffar .
jag delar även kritiken mot att inget avseende har fästs vid artikel 82 , framför allt med tanke på att vi kan tillgripa oriktiga metoder vid en koncentration av marknaden .
i egenskap av ledamot från baskien , vill jag uttala mitt fulla stöd för åtgärder som att tillämpa en vederbörlig konkurrens på marknaden .
jag vill påpeka detta om det nu skulle råda några tvivel angående den kritik vi riktat mot kommissionen i allmänhet och mot monti i synnerhet , på grund av dennes attack mot stimulansåtgärderna till de baskiska företagen och det faktum att han betraktar dessa som ett statligt stöd .
det vi skulle reagera negativt på är om kommissionen gick vidare utan att ha förstått det inre väsendet hos det generella systemet i vår ordning , med ett medansvar , som innebär att våra baskiska taxeringsnormer är av samma karaktär , att grundsatserna och målsättningen med dessa är samma som för normerna i unionens stater , och att dessa normer gäller alla skattebetalare som på ett eller annat vis omfattas av dem .
herr talman , herr kommissionär ! ja , vi behöver konkurrens !
vi behöver konkurrens för att få så låg arbetslöshet som möjlighet , för att få en välutvecklad hälsovård , social rättvisa , hög social standard , och vi behöver naturligtvis också - det är nationalekonomiska konkurrenskriterier - en företagsekonomisk konkurrens : högsta kvalitet på produkterna , samma villkor för tillgången till marknaden för alla företag , miljövänliga produkter .
det betyder att vi måste lyckas koppla samman de nationalekonomiskt erforderliga konkurrenskriterierna med de företagsekonomiska .
jag får ofta intrycket att i motsats till hur det förhöll sig i det land som jag kommer från - östtyskland - där den nationalekonomiska konkurrenskraften var närmast allenarådande och den företagsekonomiska inte beaktades , gör man nu ofta motsatsen ; samhället tänker nästan enbart företagsekonomiskt .
detta säger jag själv som företagare , som absolut är intresserad av detta .
men på det viset kan ett system inte fungera ! det måste finnas en koppling .
jag vill ge er ett exempel : europeiska unionen har med all rätt stött stålverket grönitz i brandenburg , fastän endast 700 arbetstillfällen återstår av 5 000 .
men det är konkurrenskraftiga arbetstillfällen , ty detta stålverk är nu nummer 2 bland verktygsstålstillverkarna i förbundsrepubliken tyskland .
den som nu i princip äventyrar produktionen i detta stålverk genom att kräva tillbaka det tidigare godkända stödet , äventyrar inte bara själva stålverket , utan han äventyrar i denna region en arbetsgivare som naturligtvis även små och medelstora företag är beroende av .
detta kan naturligtvis inte vara europeiska unionens konkurrenspolitik !
om vi vill ha konkurrens , då måste vi få till stånd denna koppling mellan de nationalekonomiska nödvändigheterna och de företagsekonomiska förutsättningarna .
det är också den enda chansen att bygga upp regionala ekonomiska kretslopp i de underutvecklade regionerna på detta sätt , som innebär att det finns en social trygghet för människorna och att köpkraften stärks .
därmed måste vi också ta avsevärt mycket större hänsyn till en ekonomisk politik som är inriktad på efterfrågan , än till en som är enbart utbudsinriktad .
herr talman ! inte sedan jag valdes in i detta parlament 1994 har jag sett ett betänkande med så anti-irländska känslor och övertoner som jonckheers betänkande som vi diskuterar i dag .
jag skulle vilja citera betänkandet ord för ord : &quot; det statliga stödet per capita är störst i italien , tyskland och irland .
irland är dock det land som får mest stöd om man lägger ihop det nationella stödet och gemenskapens regionala och sociala stöd . &quot;
jag anser att föredraganden bara leker med siffror .
jag har svårt att inse hur han kan stoppa in regionala och sociala fonder i denna matematiska ekvation .
jag skulle vilja påminna ledamoten om att europeiska unionen har antagit de nya riktlinjerna för regionalstöd för perioden efter år 2000 .
detta var bara en förlängning av de politiska målsättningarna att komplettera den inre marknaden i europa .
regionala skillnader måste övervinnas om den inre marknaden skall lyckas och frodas .
det faktum att ett stöd på 40 procent med ytterligare 15 procent till små och medelstora företags fasta investeringskostnader kommer att beviljas för företag som startas i mål 1-regioner i europa efter år 2000 är välkommet .
jag påminner jonckheer om att irländska företag och utländska företag i irland fortfarande måste ta sig över två hav för att komma till marknaden på det europeiska fastlandet .
ingen annan medlemsstat har ett så ogynnsamt läge .
herr talman , mina damer och herrar , kära kolleger ! kartellförbudet utgör kärnan i en fungerande konkurrensordning i europa .
det praktiska hanteringen av övervakningen av kartellförbudet har kommissionen funnit vara otillfredsställande ; det kan man till att börja med hålla med om .
men i fråga om lösningen skiljer sig åsikterna åt .
kommissionens förslag avviker formellt inte från kartellförbudet , men till sitt resultat är detta förslag en övergång från ett förbud med godkännandeförbehåll till ett godkännande med förbudsförbehåll .
detta är en växling från förbudsprincipen till missbruksprincipen .
en så graverande systemändring avvisas beslutsamt av mig och andra kolleger .
jag godtar inte att ett problem med det praktiska genomförandet skall ge anledning till att ändra rättsordningen .
vi ändrar på rätten för att det åter skall gå att verkställa den ; det anser jag inte vara godtagbart .
kommissionen avstår från sitt monopol att ge undantag för vissa slag av stöd .
mot bakgrund av detta planerade system med direkt tillämplighet av undantagsregeln är konkurrensbegränsningar utan vidare undantagna , såvida det föreligger förutsättningar enligt artikel 81.3 eg-fördraget .
nödvändigheten av anmälningar till bryssel faller bort , vilket innebär att kommissionen i denna sak kommer att flyga med autopilot i framtiden .
det finner jag inte godtagbart .
kommissionens koncept kompletteras genom en ökad kontroll i efterhand av de nationella myndigheterna och domstolarna i medlemsstaterna .
här kommer vi emellertid , om det äger rum på detta vis inom ramen för en åternationalisering , att få en konkurrenspolitisk trasmatta i europa .
jag tror inte det är godtagbart .
här försvagas en kärnpunkt i den europeiska politiken .
den av kommissionen planerade systemändringen i den europeiska kartellrätten är konkurrenspolitiskt sett synnerligen riskabel .
vi har tillräckligt med andra optioner i det befintliga systemet för att säkra öppna marknader och fri konkurrens .
för övrigt kommer kommissionen med sitt förslag åter tillbaka till gamla förslag , som lades fram redan någon gång på 50- och 60-talet .
de fick ingen majoritet .
eftersom frankrike då mycket starkt ställde undantagsregeln i förgrunden , kompenserades man av eftergifter inom jordbrukspolitiken .
fyrtio år senare dyker detta förslag nu upp igen , och det kommer - det är jag säker på - att ge utrymme för kartellbildningar till nackdel för konsumenterna i europa .
jag anser inte att det är godtagbart !
herr talman , kära kolleger ! i denna viktiga konkurrensdebatt vill jag i dag mera särskilt uttala mig om langens text , om gemenskapens regler för stöd till stålindustrin .
stålsektorn är särskilt känslig för konkurrensstörningar , något som eg-domstolen erkände år 1996 .
jag drog för övrigt själv samma slutsats för några år sedan , i ett betänkande om den europeiska stålindustrins styrka och svaghet .
det var därför berättigat att inrätta ett stödsystem för denna sektor , i syfte att garantera de livskraftiga företagens överlevnad , även om det stod i strid med artikel 4 i eksg-fördraget .
detta är syftet med den sjätte regeln för stöd till stålindustrin . men samtidigt är det viktigt att förhindra att konkurrensvillkoren kränks och att marknaden utsätts för allvarliga störningar , därav vikten av att fastställa regler för den här typen av stöd .
det är således nödvändigt att även i fortsättningen begränsa statsstöden till följande områden : forskning , utveckling , miljöskydd samt nedläggningar av företag .
av samma skäl är det ytterst viktigt att medlemsstaterna uppfyller förpliktelsen att till kommissionen anmäla de stöd som de beviljar sina stålföretag .
kommissionen föreslår snävare tidsramar .
jag instämmer i det förslaget .
i likhet med föredraganden gläder jag mig åt kommissionens rapport , men beklagar ändå att den inte täcker alla aspekter av dessa stöd .
trots att gemenskapens regler om stöd till stålindustrin formuleras på ett mycket tydligt sätt , har kommissionen beviljat stöd till stålföretag som inte tillhör någon av de kategorier som åsyftas i reglerna .
med omsorg om rättvisa bör man antingen tillämpa reglerna eller ändra på dem .
för att till sist avsluta , herr talman , krävs det en översyn av reglerna innan eksg-fördraget löper ut , för jag anser att stödsystemet bör finnas kvar efter år 2002 . jag är följaktligen positiv till att en förordning från rådet skall erbjuda en garanti i det avseendet .
därför väntar vi - jag inväntar förslag från europeiska kommissionen med den innebörden .
herr talman ! även jag kommer att tala om langens betänkande beträffande stödet till stålindustrin .
jag håller med föredraganden på två punkter .
för det första vad gäller behovet av att garantera lika villkor för stödet till alla medlemsstater , och för det andra vad gäller stödets genomblickbarhet .
vi kritiserar , precis som föredraganden , att kommissionen trots de normer som härrör sig från det sjätte regelverket om stöd till stålindustrin , vid flera tillfällen har beviljat stöd till företag som inte överensstämmer med kategorierna för reglerna .
hur som helst , herr talman , det som mest bekymrar oss är sänkningen av priserna med 30 procent till följd av importen .
orsaken till denna prissänkning är den illojala konkurrensen från sydkorea och taiwan inom stålindustrin , på grund av andra villkor för arbete och stöd .
orderingången inom stålindustrin och sjöfartssektorn - den frågan diskuterade vi nyligen - har minskat drastiskt med en minskad sysselsättning som följd .
jag bor i en region där sjöfartssektorn för närvarande lider av stora problem : asturien .
för marknader med internationell räckvidd bör det finnas arbetsnormer med internationell räckvidd och stöd med internationell räckvidd .
jag vet att det är svårt att åstadkomma något sådant nu , men om vi inte lyckas åstadkomma rättvisa arbetsnormer för alla arbetstagare , både här och i övriga världen , om vi inte kan åstadkomma ett rättvist stöd för alla länder , både här och i övriga världen , kommer det att bli mycket svårt att bibehålla sysselsättningen , både i europa och i övriga världen .
herr talman , herr kommissionär , herr generaldirektör , mina damer och herrar ! jag vill framför allt konstatera följande beträffande von wogaus betänkande : jag välkomnar kommissionens ansträngningar att utan något tabu inleda en diskussionsprocess om de hittills benhårda reglerna om förfarandena , och föreslå konkreta reformåtgärder .
jag gratulerar föredraganden karl von wogau , som tar itu med saken , men också helt konkret kräver klargöranden , hänvisar till erforderliga åtföljande åtgärder och kritiskt kallar de aktuella uttalade problemen vid deras rätta namn .
vitboken och betänkandet bidrar i inledningsskedet till en process av nödvändig eftertanke , nödvändiga diskussioner och reformer , som ännu inte är avslutad , eftersom somliga frågor fortfarande måste redas ut av oss , av domarna , medlemsstaterna och framför allt av de berörda små och medelstora företagen .
konkurrenspolitiken måste även i fortsättningen hanteras centralt och kommer inte att åternationaliseras , eftersom detta skulle äventyra den inre marknaden och handelsplatsen europa i den globala världsekonomin .
men den måste europeiseras på ett sätt som motsvarar subsidiariteten .
jag välkomnar därför också att ansvaret läggs på den enskilde , utan att kommissionen undandrar sig sitt ansvar .
erfarenheterna i praktiken - endast 9 fall avvisades , och 94 procent av de fall som kommissionen skulle bearbeta klarades av inte formellt , utan endast med hjälp av icke offentliggjorda , rättsligt icke bindande administrativa skrivelser eller helt enkelt på grund av att tiden gick - visar tydligt att man måste sätta tidsmässiga , personella och finansiella gränser för kommissionens arbete i en tidsålder av globalisering och eu-utvidgning .
avslutningsvis vill jag säga vad jag förväntar mig av denna reform : en rättvis konkurrens och lika konkurrensvillkor , rättssäkerhet för alla företag , en enhetlig tillämpning av konkurrenspolitiken , förenklade förfaranden enligt principen one-stop-shop , en samordning av de nationella och för mig oberoende konkurrensmyndigheterna , ett nära samarbete mellan de nationella myndigheterna och domstolarna och kommissionen , liksom en klar ansvarsfördelning mellan nationella myndigheter och domstolar vid tillämpningen av den europeiska konkurrens- och kartellrätten ; av kommissionen förväntar jag mig att den koncentrerar sig på väsentligheterna genom att fullgöra sina uppgifter som högsta väktare av den europeiska konkurrenspolitiken .
jag väntar med spänning på att få se hur diskussionerna , som förs på bred basis , kommer att mynna ut i det första lagförslaget .
kommissionens rapport bekräftar att de statliga företagsstöden ökar , tyskland undantaget .
men det enda som oroar kommissionen är konkurrensvillkoren .
vi sätter oss däremot in i arbetarklassens intressen .
samhället tjänar ingenting på de enorma överföringarna av offentliga medel till privata företag .
titta på bilbranschen ; där har statliga subventioner och olika former av statsstöd ökat med 24 procent under den granskade perioden .
av vilka skäl då ?
inte för att bevara arbetstillfällen .
alla dessa företag har avvecklat arbetstillfällen , ja t.o.m. avskedat folk .
och det är inte för att förbättra arbetsvillkoren , för arbetsvillkoren försämras när färre arbetare skall producera mer .
var dessa företag i behov av statliga stöd för att överleva ?
nej , biltillverkarna håvar in kolossala vinster sedan flera år tillbaka .
de statliga stöden får inte endast negativa bieffekter då de främjar en jakt på subventioner genom omlokaliseringar från ett land till ett annat , vilket medges i jonckheerbetänkandet ; de är också oacceptabla eftersom de innebär att offentliga medel används för att berika en handfull privata aktieägare .
eftersom man överallt gynnar de rikaste med hjälp av statens pengar , inskränker man också det sociala skyddet överallt i europa - man överger den offentliga sektorn , man lägger ner sjukhus .
genom att rösta emot jonckheerbetänkandet vill jag hävda att det krävs en annan politik , dvs. att alla stöd till privata företag stoppas och att de därmed frigjorda pengarna används för att utveckla tjänster av allmänt intresse och för att anställa personal inom den offentliga sektorn .
herr talman ! dagens debatt är utomordentligt viktig , för konkurrensprincipen har förmodligen varit hörnstenen för den inre marknaden .
som ett sätt att tillämpa konkurrensprincipen har man utformat artiklarna 85 till 94 , konkurrenspolitiken närmare bestämt , granskningar av sådant statligt stöd och sådana skattebestämmelser som skulle kunna förändra konkurrensen .
till en början de indirekta skattebestämmelserna ; och nyligen , tack vare kommissionär monti , de direkta bestämmelserna , och då i synnerhet uppförandekoden .
detta har fungerat tämligen väl , men tiden går , precis som i den välkända filmen casablanca , och det är nödvändigt att anpassa de bestämmelser som vi hittills har tillämpat till de nya omständigheterna .
jag har lagt märke till en stark enighet på den punkten i alla anföranden .
för det första är det nödvändigt att man i utformningen av bestämmelserna gör upp tydliga och heltäckande regler .
förmodligen är förekomsten av oklara regler , oreglerade områden eller regler som endast fastslår vaga juridiska begrepp allvarligare i denna del av bestämmelserna än i andra delar .
inte minst - så som fallet är i reformens andra del - då tillämpningen av bestämmelserna överlåts åt de nationella myndigheterna .
för det tredje , anser jag att kommissionen har en viktig roll att fylla i och med att man motstår frestelsen att inrätta oberoende byråer , något som skulle förändra kommissionens innersta väsen , som ett sätt att garantera en enhetlig tillämpning från de internationella organens sida .
och slutligen för det fjärde- och det har redan påtalats - har den internationella rättsordningen förändrats .
det kunde vi se i och med den misslyckade konferensen i seattle och nu ser vi det i samband med de bilatera konferenserna för olika regioner eller länder .
konkurrensprincipen bör ha en universell tillämpning .
och vi bör se till att miljönormerna , arbetsnormerna följs , för att undvika dumpning på det området , att rätten till egendom respekteras fullt ut , att det sker en granskning av det statliga stöd som - precis som det har sagts här - snedvrider konkurrensen inom flera sektorer och förstör sysselsättningen på hemmaplan , och vi bör definitivt se till att snarlika villkor tillämpas som förhindrar att stödåtgärder , snedvridningar på den inre marknaden i andra länder sprids till internationell nivå genom fusk .
herr talman , herr kommissionär monti ! jonckheers betänkande om statliga stöd till tillverkningsindustrin och vissa andra sektorer innehåller mycket gott .
för det första framhåller man i betänkandet parlamentets fasta ståndpunkt att de statliga stöden målmedvetet måste minskas för att den inre marknaden skall kunna fungera korrekt .
många av betänkandets slutsatser vållar dock åtminstone inom vår grupp allvarlig oro .
att sådana här översikter är nödvändiga bevisas till exempel av det faktum att mängden av och nivån på det statliga stödet per capita varierar kraftigt mellan olika medlemsstater .
stöd som väller fram till följd av nationella egoistiska utgångspunkter ger företagen orättvisa fördelar , snedvrider på det sättet konkurrensen och leder till en ineffektiv och oekonomisk fördelning av de knappa europeiska resurserna .
det är inte heller helt oväsentligt vilka typer av stöd det handlar om .
statliga stöd som förutsätter egna ansträngningar av stödmottagaren måste prioriteras .
de statliga garantierna till exempel , angående vilka kommissionen nyligen offentliggjort ett ställningstagande , måste naturligtvis räknas till de statliga stöden men är enligt min mening ett bättre alternativ än direkta bidrag till företag .
rapporten om konkurrenspolitiken framhäver vidare kommissionens tro på kraftig reglering i stället för att betona de ekonomiska effektivitetsargument som påverkar konkurrenskraften .
den europeiska ekonomin kommer aldrig att uppnå önskad konkurrenskraft om vi inte visar att vi litar på marknadens funktion .
om konkurrenspolitiken skall underordnas social- och miljöpolitiska ambitioner kan vi bara drömma om verklig effektivitet och ekonomisk tillväxt .
konkurrenspolitiken måste också ses som en del av den ekonomiska helheten och den måste bedömas bland annat i förhållande till handelspolitik och immateriella rättigheter . man kan inte enbart betona dess sociala dimension .
socialpolitiska mål uppnås bäst genom en kraftigare ekonomisk tillväxt , inte genom att kompromissa om konkurrenspolitiska lösningar .
i rapkays betänkande betonas också konkurrensrättens internationella dimension .
jag tycker också att det är bra om man på internationell nivå uppnår samförstånd när det gäller vissa konkurrensrättsliga kärnprinciper .
om man däremot strävar efter enhetliga miniminormer leder detta lätt till att man går den enklaste vägen och väljer den minsta gemensamma nämnaren , vilket urvattnar alla konkurrenspolitiska mål .
herr talman , kommissionär monti ! uppdateringen av konkurrensreglerna borde vara en viktig uppgift för europeiska unionen , inte bara mot bakgrund av och som en konsekvens av de förändringar som inträffat genom åren , utan också med tanke på unionens förestående utvidgning .
jag tackar föredraganden karl von wogau för det engagemang han lagt ner och jag uppskattar verkligen hans resonemang .
jag vill också uttrycka min uppskattning för de synpunkter som jag har fått från professor tesauro , ordförande för den italienska myndigheten , och som jag är övertygad om att professor monti i en anda av samförstånd kommer att ta vederbörlig hänsyn till .
det problem vi står inför är utan tvekan hur vi skall kunna ytterligare avreglera marknaden och framför allt se till att de olika nationella marknaderna blir homogena , de marknader som för tillfället uppvisar stora skillnader , skillnader som tydligt framkommer om man jämför den engelska marknaden med den italienska och franska .
på den senare finns det starka inslag av statlig protektionism , något som inte finns på den engelska och som är ytterligt begränsat i italien .
ett annat problem är ekonomierna i de länder som berörs av utvidgningen , som riskerar att för evigt bli subventionerade ekonomier om det inte kan ske en gradvis anpassning .
enligt min mening är det även nödvändigt att skapa en nivå där man skall införa två viktiga inslag som karakteriserar vårt ekonomiska system : de små och medelstora företagen , som utgör det sammanbindande elementet i den europeiska ekonomiska verkligheten , och det sociala skydd som europa alltid har garanterat de ekonomiskt svagaste grupperna .
skyddet av marknadens sociala dimension utgör hela skillnaden mellan en total marknadsliberalism och ett system som skall kunna förbättra människors livskvalitet .
en aspekt som måste beaktas i det nya regelverket utgörs av ekonomierna i de ultraperifera regionerna och i öregionerna , som behöver skyddas .
därför tror jag att det skulle vara lämpligt att även tänka på att skapa två fokus för den externa marknaden och att inleda ett givande samarbete med ryssland och medelhavsländerna , just för att de ekonomierna skall bli mindre perifera .
jag hoppas - och i det sammanhanget vill jag tacka professor monti - att man i det nya regelverket ägnar ett så stort utrymme som möjligt åt den ekonomiska politiken och att man verkligen garanterar dess sociala funktion .
herr talman ! konkurrens är hjärtat och kraften i den europeiska politiken för den inre marknaden .
en fri öppen marknad kan bara existera under konkurrensens överhöghet , begränsad av tydliga , enhetliga spelregler .
karl von wogau förordar detta på ett mycket bra sätt i sitt betänkande .
men europa förändras .
ekonomierna växer , vi expanderar till 25 till 30 medlemsstarter .
europeiska kommissionen kommer att bli överbelastad om den nuvarande politiken skall fortsätta .
det är därför nödvändigt med en modernisering av konkurrenspolitiken .
det råder ingen diskussion om detta .
men trots detta kan jag ändå inte släppa en oro i fråga om den planerade decentraliseringen .
på vilket sätt kommer kommissionen som fördragens väktare att garantera att man på ett enhetligt sätt fattar beslut i konkurrensärenden i london , palermo , helsingfors och inom kort i budapest och ankara ?
det är nödvändigt att förhindra olikhet inför lagen , annars skulle en strid ström av konkurrensmål gå till den domstol där den mildaste bedömningen görs .
det räcker inte med att säga att medlemsstaterna redan har 40 års erfarenhet .
i nederländerna ligger konkurrensmyndigheten fortfarande i sin linda .
detta land har att göra med en mycket liten marknad som tyvärr ofta samtidigt definieras som den relevanta marknaden .
detta i motsats till tyskland , där en mycket erfaren kartellamt utövar sina befogenheter på en gigantisk marknad .
europeiska kommissionens tilltro till att tolkningen av lagstiftningen kommer att vara lika i alla väderstreck är vad vi i katolska kretsar kallar &quot; övermodigt förtroende &quot; , och det är förbjudet .
det krävs mer arbete för att uppnå enhetlighet .
jag tänker på specialiserade , nationella domstolar med möjlighet att överklaga direkt till en särskild konkurrensdomstol vid eg-domstolen .
denna särskilda domstol behövs på grund av att det är nödvändigt att bygga upp en bred expertis .
dessutom tillåter inte de mycket stora ekonomiska och sociala intressen som hör samman med ärenden av den arten att ett domslut låter vänta på sig i två år , vilket nu är helt normalt .
vad anser kommissionären om detta ?
jag vill avsluta med en viktig punkt för det lilla och medelstora företaget .
för att skapa trygghet för det lilla och medelstora företaget bör europeiska kommissionen själv utarbeta en undantagsförordning för det lilla och medelstora företaget i syfte att också möjliggöra horisontala undantag vid sidan av vertikala .
småföretagare måste genom samarbete kunna försvara sig mot de stora kedjorna .
syftet med den europeiska konkurrenspolitiken kan inte vara att göra livet omöjligt för småföretag .
vad småföretag beträffar bör man dessutom begrunda om det inte skulle kunna vara lättare att hantera ett system med en varning i förväg , gult kort , i stället för att omedelbart ge ett rött kort som kommer att fungera som böter och hota företagets fortlevnad .
herr talman ! i egenskap av sista talare har jag privilegiet , herr kommissionär , att få tala om att majoriteten av den här församlingen stöder ert initiativ och har visat ett fullständigt , och jag tror även högst berättigat förtroende för er som kapten på den här skutan .
men vi vill utgöra besättningen på skutan , eftersom vi befinner oss på samma skuta som ni .
därför anser jag att en interinstitutionell dialog är oumbärlig , så att vi kan precisera och nyansera denna så viktiga reform och föra den i hamn .
de förslag som har lagts fram här kan delas in i tre stora grupper .
i första gruppen finns den oro som vissa av oss har gett uttryck för , och då i synnerhet randzio-plath , ordförande i utskottet för ekonomi och valutafrågor , en oro för att detta nya system som ett rättsligt undantag inte skall överensstämma med fördraget .
jag delar hennes oro och anser att den saken bör undersökas .
i andra gruppen ingår frågan om företagens rättssäkerhet .
det är sant , herr kommissionär , att kommissionen inte är en maskin som tillverkar rättssäkerhet .
det kan vi alla vara överens om .
men det är likaså sant - och det har alla sektorer i den här församlingen upprepat - att den europeiska industriella vävnaden är en vävnad som består av små och medelstora företag , och att kommissionen många gånger är den som företräder auctoritas , legitimering , legitimitet , av det som är den inre marknaden .
på den punkten vill jag framföra min åsikt om något karas sade .
det har endast förekommit nio beslut om avslag .
där har jag nytta av min erfarenhet som advokat .
hur många gånger har det inte hänt att en advokat med två bolag och ett projekt har ändrat projektet efter en orientering ex ante från kommissionens sida , för att det skall överensstämma med konkurrensbestämmelserna !
det är därför en aspekt att ta hänsyn till .
i den tredje gruppen ingår problemet med en enhetlig tillämpning av gemenskapsrätten .
thyssens utmärkta inlägg kunde knappast ha varit bättre .
jag anser att det är bra med ett biologiskt mångfald , och även med ett kulturellt mångfald , däremot inte med ett mångfaldigt tillämpande av rätten , av det som är själva kärnan i den inre marknaden , det vill säga , konkurrensbestämmelserna .
där krävs en närmare precisering .
endast i vissa länder , som i tyskland , har man en specialiserad rättsskipning .
måhända är det en lösning som är värd att undersöka , men vi bör även undersöka andra möjligheter .
det vi inte får göra , herr kommissionär - och med detta vill jag avrunda - är att ge så mycket som ett lillfinger , och än mindre räcka vapen åt dem som talar om de europeiska institutionerna som en fråga för de mäktiga , för de inflytelserika , för de rika , och inte för den enskilda medborgaren , inte för de små och mellanstora företagen , som skulle känna sig utelämnade åt sina värsta föreställningar- som aldrig kommer att förverkligas , för de rätta åtgärderna kommer att vidtas för att undvika något sådant - till domstolar som avkunnar olika domar , mycket sent , utan några realistiska möjligheter till kontroll annat än med det som fransmännen kallar le parcours du combattant , det vill säga efter jag vet inte hur många år , när domstolen i luxemburg uttalar sig , en domstol som vi alla vet för närvarande är starkt överbelastad .
herr kommissionär , vi står inför en reform som jag inte nog kan poängtera vikten av .
effekten av denna reform sprider sig till konkurrensen , den sprider sig till sammanhållningen på den inre marknaden , jag tror att den på djupet påverkar det som är meningen med den europeiska integrationen , meningen med den europeiska integrationens legitimitet .
därför , herr kommissionär , räknar vi med denna interinstitutionella dialog som ett sätt att närmare precisera en reform som vi alla hoppas och tror att vi kommer att ro i hamn med er som kapten och oss som besättning .
herr talman , ärade ledamöter ! låt mig varmt tacka utskottet för ekonomi och valutafrågor och hela europaparlamentet för det stora intresse de visar för konkurrensfrågorna .
denna gemensamma debatt är , herr talman , enligt min åsikt ett levande och starkt bevis på detta .
vi har lyssnat på resonemang av stor djupsinnighet som samtidigt har rört ekonomisk politisk filosofi och institutionernas arbete .
vår gemensamma avsikt är att uppdatera , förstärka konkurrenspolitiken , grundbulten i den sociala marknadsekonomin och det europeiska konstruktionsarbetet .
den röda tråden i arbetet med att reformera konkurrenspolitiken , som vi skall genomföra gemensamt , är syftet att garantera ett säkrare skydd för konkurrensen , minska den byråkratiska börda som tynger företagen , och att föra beslutsprocesserna närmare medborgarna .
jag vill personligen varmt tacka von wogau för det engagemang han visat i arbetet med vitboken och för den goda kvaliteten i hans betänkande .
låt mig sammanfatta de synpunkter som framförts i debatten om von wogaus betänkande i fyra punkter , som jag inte anser vara kritik mot kommissionen , utan snarare som bidrag av avgörande betydelse , eftersom det finns invändningar som det är viktigt att framföra och som vi tillsammans vill reda ut : frågan om effektiviteten , frågan om risken för åternationalisering , frågan om en enhetlig tillämpning , frågan om rättssäkerheten .
låt mig som hastigast gå igenom dem en efter en .
effektiviteten : jag är övertygad om att denna reform kommer att göra det möjligt för oss att förstärka , snarare än försvaga , konkurrensskyddet inom ramen för den inre marknaden .
det nuvarande anmälningssystemet , ärade parlamentsledamöter , tillåter oss inte längre att uppnå det målet eftersom det inte garanterar information till kommissionen om de allvarligaste restriktionerna - låt mig påminna om att under trettiofem år har endast nio beslut om förbud fattas som en följd av en anmälan och där det har saknats en stämning - inte garanterar öppenhet och inte medför en reell rättssäkerhet för företagen som , i de flesta fall , mottar ett enkelt administrativt meddelande som sedan arkiveras .
det system som föreslås gör det möjligt att förbättra konkurrensskyddet , framför allt därför att det kommer att tillåta kommissionen att koncentrera sin uppmärksamhet på de allvarligare inskränkningarna , just därför att det i högre grad kommer att engagera de nationella konkurrensverken i arbetet att hålla nere kränkningarna och , slutligen , för att det gör det möjligt för dem som drabbas av kränkningarna att vända sig direkt till de nationella rättsinstanserna , vilkas uppgift det är att skydda de enskildas rättigheter .
frågan om åternationaliseringen : först av allt , även om det skulle vara överflödigt , skulle jag vilja påminna om och understryka , tre gånger om det är möjligt , att vitboken inte i något avseende berör frågan om koncentrationer och statliga stöd - vi överväger inte en tillbakagång i det avseendet - utan , när det gäller förordning 17 , så finns det en risk för åternationalisering .
ni kan föreställa er att vi naturligtvis har ställt oss den här frågan : vi har ställt oss frågan och vi följer den uppmärksamt , även tack vare den oro som ni har givit uttryck för .
men jag tror uppriktigt sagt inte att denna oro är berättigad .
kommissionens förslag ger kommissionen en central roll när det gäller att bestämma konkurrenspolitikens inriktning .
reformen innebär ingen minskning i kommissionens verksamhet , utan en koncentration av uppmärksamheten till de viktigaste fallen .
reformen kommer att leda till en gradvis utveckling låt mig understryka detta för jag tyckte om den formulering som användes av ordföranden randzio-plath och som jag för övrigt helt instämmer i - av en europeisk konkurrenspolitik .
reformen kommer att leda till en överföring , en omplantering på den europeiska konkurrenskulturens mark - där det i dag växer diverse olika plantor , som verkligen inte är enhetliga - av de olika nationella konkurrenskulturerna .
det kommer att leda till att man gradvis överger de femton olika nationella rättssystemen till förmån för en vidare tillämpning av gemenskapsrätten , som kommer att kunna tillämpas av allt fler aktörer .
detta , tillåt mig understryka det , är att göra konkurrensrätten gemensam , och inte att åternationalisera den .
frågan om den enhetliga tillämpningen : vi skall vara medvetna om risken för en icke enhetlig tillämpning av konkurrensreglerna , men jag tror samtidigt att den risken inte skall överdrivas .
i likhet med flera andra föreskrifter i fördraget , artikel 81.1 och 82 , tillämpas de trots allt sedan decennier av nationella myndigheter och domare , och jag tycker inte att detta har skapat några större problem .
inom ett överreglerat område är en enhetlig tillämpning i första hand beroende av graden av klarhet i de grundläggande rättsreglerna .
kommissionen kommer att anstränga sig för att verkligen precisera den rättsliga ramen , såväl via allmänna åtgärder som i de praktiska besluten .
för det andra måste vi få till stånd effektiva konfliktförebyggande mekanismer och här föreslås i vitboken system för information och samråd .
låt mig i det sammanhanget säga ett ord om den i mitt tycke utmärkta idé som framförts av riis-jørgensen och huhne , dvs. idén om tillämpningsövervakning - monitoring of the implementation .
så detta är vad idén att övervaka verkställandet går ut på .
jag måste säga att jag tycker att det är en mycket god idé som vi troligen kommer att ta upp .
även om vi har stor respekt för de nationella konkurrensmyndigheternas arbete och så vidare är det uppenbart att vi kommer att syna hur eg : s lagar tillämpas av nationella myndigheter och domstolar mycket noggrant .
det är därför kommissionen vill ha kvar rätten att dra tillbaka ett fall från en nationell konkurrensmyndighet vid eventuell felaktig tillämpning .
detta borde minska er oro i någon mån , fru peijs .
( en ) vad beträffar evans fråga om konsekvenserna för företagen är det viktigt att den samhällsekonomiska kostnads-intäktsanalysen genomförs på ett seriöst sätt .
syftet med att ge ut en vitbok är när allt kommer omkring att inhämta synpunkter från företag lika väl som från andra källor .
vi har fått in många utmärkta påpekanden och bidrag som ger oss underlag för att göra en kostnads-nytto-analys för industrin .
vi kommer att gå igenom allt detta material noggrant innan vi lägger fram ett förslag till ny lagstiftning .
det finns en aspekt av konsekvenserna för företagen som är mycket viktig .
denna togs upp av thyssen , peijs och palacio vallelersundi : frågan om små och medelstora företag .
många talare har betonat detta .
kommissionen är särskilt uppmärksam på de små och medelstora företagens rättssäkerhet .
vi föreslår ett system som stärker de små och medelstora företagens rättssäkerhet betydligt .
är detta enbart en politisk gest ?
i systemet föreslår vi att våra grundläggande regler ändras på ett sådant sätt att de flesta små och medelstora företag kommer att omfattas av generella undantag , såsom vad beträffar de vertikala begränsningarna .
de flesta små och medelstora företag har faktiskt en marknadsandel på mindre än 30 procent .
vi har en de minimis-notis där vi förklarar att eftersom små och medelstora företag inte är involverade i marknadsdominans omfattas de normalt inte av det stränga förbudet i artikel 81.1 .
vi arbetar på ytterligare generella dispenser och riktlinjer som alla kommer att ta hänsyn till de små och medelstora företagens speciella situation , och vår vitbok om modernisering kommer också att förbättra för de små och medelstora företagen genom att för det första den byråkrati det nuvarande anmälningssystemet ger upphov till försvinner och för det andra genom att artikel 81.3 blir direkt tillämplig , vilket kommer att gynna speciellt de små och medelstora företagen .
( it ) den fjärde frågan gäller rättssäkerheten .
naturligtvis , evans , är rättssäkerheten - jag är den förste att hålla med om det - viktig för företagen , inte bara för juristerna som även spelar en mycket viktig roll i det europeiska konstruktionsarbetet .
rättssäkerheten är viktig för företagen : detta är en fråga som ordföranden för utskottet för rättsliga frågor och den inre marknaden , palacio vallelersundi som jag vill tacka för att hon alltid behandlar frågorna som rör den inre marknaden på ett uttömmande vis , dvs. i detta fallet inklusive konkurrensfrågan - även i sitt senaste inlägg underströk betydelsen av .
jag är övertygad om att detta förslag kommer att öka företagens rättssäkerhet , och detta av tre anledningar : det gör det möjligt att utan ett föregående beslut godkänna samtliga konkurrensbegränsande avtal som uppfyller villkoren om utvidgning , tack vare den direkta effekten av artikel 81.3 ; det skapar möjligheter att hjälpa företagen om det uppkommer tolkningsproblem , genom publicering av motiverade beslut ; det kommer att åtföljas av undantagsbestämmelser och riktlinjer i avsikt att förtydliga reglerna och garantera deras säkerhet .
( fr ) thyssen nämnde också frågan om företagsjuristernas legala privilegium .
låt mig endast erinra om att eg-domstolen avgjorde den frågan 1982 , det vet ni bättre än jag . denna rättspraxis är fortfarande giltig och det finns ingenting som gör det motiverat att ifrågasätta den .
enligt vitboken skall frågan åter granskas med avseende på en aspekt : utbyte av sekretessbelagd information .
vilka garantier företagen bör få är för närvarande föremål för diskussioner .
( it ) herr talman ! jag kommer så till rapkays betänkande och jag vill först tacka ledamot rapkay för kvaliteten i arbetet och för det stöd som ges kommissionens 28 : e årsrapport om konkurrenspolitiken .
jag tycker mig finna en betydande samsyn , men i rapkaybetänkandet understryks vissa saker som det är vår skyldighet att beakta mycket noga .
jag vill av tidsskäl här endast peka på två : den ena gäller en ytterligare ökning av öppenheten .
detta parlament vet att vi alla anser att öppenheten är en mycket viktig fråga inom konkurrenspolitiken , och jag personligen har från första början hävdat detta , alltsedan den 1 september , dvs. den första dagen av min utfrågning inför utskottet för ekonomi och valutafrågor .
när det gäller konkurrenspolitikens internationella dimension kan jag bekräfta för er , ledamot rapkay , att kommissionen är beredd att lägga fram en rapport i frågan för parlamentet , denna fråga som även randzio-plath har pekat på och inom ramen för vilken jag kan nämna att vi har upprättat mycket tillfredsställande bilaterala kontakter med motsvarande myndigheter i usa , kanada , japan och vi kommer att arbeta för att världshandelsorganisationen skall anta konkreta regler på konkurrensområdet .
jag vill lika varmt tacka er , ledamot jonckheer , för ert betänkande om sjunde översikten över statligt stöd i europeiska unionen inom tillverkningsindustrin och vissa andra sektorer .
jag tänker inte här gå in på frågan om medbeslutande , men det beror inte på att jag inte anser den viktig .
den frågan har en institutionell betydelse som naturligtvis går utöver frågan om konkurrensen . jag har med andra ord inte rätt att uttala mig i en fråga som naturligt hör hemma inom ramen för regeringskonferensen .
när det gäller era förslag , ledamot jonckheer , så vet ni redan att mina avdelningar - även om det sker med de alldeles för små , men mycket kvalificerade personalresurser de förfogar över - arbetar aktivt med att ta fram ett register över de statliga stöden och ett poängsystem över statliga stöd .
jag väntar också med spänning på resultatet av den åttonde översikten , som har följande etapper : den sammanställs av tjänstemännen nu , i januari , och antagande av kommissionen i mars 2000 , för att se om de senaste tendenserna bekräftas .
jonckheer , thyssen och gemelli har nämnt kandidatländernas förberedelser inom området konkurrens och när det gäller de statliga stöden .
låt mig bara helt kort säga att vi arbetar med dem mycket aktivt och konkret : kandidatländerna förbereder sig , de har redan infört samtliga lagar på konkurrensområdet och de håller på att inrätta respektive myndigheter .
jag kan också nämna , när det gäller oron - som jag , som ni vet , delar - för energin och framför allt miljön , att vi håller på att avsluta arbetet med att revidera lagstiftningen när det gäller statligt stöd på miljöområdet .
jag vill också understryka , när det gäller problemen med statliga stöd , den punkt som togs upp av bland andra riis-jørgensen , om ersättning för juridisk hjälp .
i april 1999 antog kommissionen en ny förordning om specifika regler för sådan ersättning .
ni kommer snart att märka - detta kan jag garantera er - att vi verkligen kommer att tillämpa de reglerna .
slutligen , herr talman , ett par ord för att varmt tacka ledamot langen för hans betänkande , som är mer sektorsinriktat , men som är lika viktigt för diskussionen .
jag kan säga att kommissionens rapport i frågan om de statliga stöden till metallindustrin , som bekant , inte omfattar de individuella beslut som fattats när det gäller undantagsförfarandet , som anges i artikel 95 i fördraget om europeiska kol- och stålgemenskapen , eftersom det rör sig om beslut som hamnar utanför tillämpningsområdet för lagen om stöd till stålindustrin .
när det gäller de kommande åtgärderna avseende stödåtgärder inom järn- och stålindustrin , som träder i kraft från och med juli 2002 , kommer vi att kräva att man fortsätter tillämpa stränga regler , vilket är ett behov som även branschen själv verkar instämma i .
när vi har lagt fram vårt förslag i frågan om nya regler och när vi har valt den juridiska form som är lämpligast , så skall det bli mig en glädje att få presentera vår vision för er .
och det , herr talman , som jag tar med mig hem efter denna debatt , en debatt som jag vill tacka parlamentet för , är ett förbehållslöst intellektuellt och politiskt stöd från europaparlamentets sida för en konkurrenspolitik , en grundläggande uppskattning för det arbete som kommissionen utför och ett förtroende för att det arbetet kan fortsätta i framtiden , saker som jag är särskilt tacksam för .
vi kommer att fortsätta , framför allt med utskottet för ekonomi och valutafrågor , men även generellt sett med parlamentet , att föra den interinstitutionella dialog som har inletts .
i det sammanhanget gladde mig er kommentar , palacio : vi måste alla ro , och helst i samma riktning .
konkurrensen är inte ett mål , som mycket riktigt rapkay har påpekat , utan ett mycket viktigt instrument i vårt europeiska konstruktionsarbete .
som von wogau sade i början på debatten , är konkurrensen trots allt inte något abstrakt : den ligger i medborgarnas intresse , den utgör en grund för den sociala marknadsekonomin .
låt mig också tillägga att i det europeiska konstruktionsarbetet har konkurrensen haft , och kommer att fortsätta att ha , ett samhällsvärde och inte bara ett ekonomiskt värde .
tack , kommissionär monti .
straffrättsliga bestämmelser till skydd för unionens ekonomiska intressen
nästa punkt på föredragningslistan är betänkande ( a5-0002 / 2000 ) av theato för budgetkontrollutskottet innehållande parlamentets rekommendationer till kommissionen om inrättande av straffrättsliga bestämmelser till skydd för unionens ekonomiska intressen .
herr talman ! jag är glad över att få ta del i debatten om detta betänkande och vill framföra mina gratulationer till theato .
jag anser att detta är ett betänkande , där samarbetet mellan utskotten har fungerat väl , och det resultat som vi i dag har fått ta del av , är ett nyktert och sansat betänkande om en synnerligen känslig fråga .
ett nyktert och sansat angreppssätt är särskilt nödvändigt vad beträffar artikel 280.4 .
för om vi ville ge ett pris åt den artikel som är mest svårbegriplig , otydlig och oklar - eller vad man nu vill kalla det - så skulle konkurrensen garanterat vara mycket jämn , för fördraget består av en brokig samling komplicerade artiklar , men denna är utan tvekan en av de starkaste kandidaterna till ett sådant pris .
samtidigt är det en synnerligen känslig fråga , eftersom det handlar om skyddet av gemenskapens ekonomiska intressen , så som theato så riktigt uttrycker det .
vi är alla medvetna om behovet - och parlamentet har tagit upp eller fört fram det problemet - av att skydda gemenskapens ekonomiska intressen .
men se upp , som fransmännen säger , &quot; ne jettons pas le bébé avec l &apos; eau du bain &quot; , det vill säga , i skyddet av gemenskapens ekonomiska intressen måste man å ena sidan respektera - och det påpekar theato - de nationella staternas behörighet , men även andra saker som påverkar medborgarna , sådant som påverkar de grundläggande garantierna .
slutsatserna i theatos betänkande värnar om dessa .
därför hoppas jag i egenskap av ordförande för utskottet för rättsliga frågor och den inre marknaden , och givetvis även som ledamot , att parlamentet i morgon antar betänkandet med stor majoritet och att kommissionen verkställer det på bästa sätt .
herr talman ! som theato sade är detta ett kritiskt betänkande .
det är ett betänkande som har föreslagits av budgetkontrollutskottet och det är ett initiativbetänkande .
en av anledningarna till att vi var mycket angelägna om att lägga fram detta var att europeiska unionen , vare sig vi tycker om det eller inte , är beryktad för bedrägerier och misskötsel .
detta är ibland överdrivet men så är det .
vi måste göra någonting åt det .
en del av medlemsstaterna har inte åtföljt vissa av de åtgärder vi har vidtagit tidigare - och låt oss inte glömma att medlemsstaterna svarar för verkställandet av omkring 80 procent av eu-budgeten .
många av dem har inte undertecknat , eller inte ratificerat konventionen om skyddet av ekonomiska intressen , och därför stod det klart att något mer radikalt behövde göras .
vi måste ta detta ansvar på allvar .
vi måste kunna åtala människor som begår bedrägerier gentemot europeiska unionen .
frågan är : vem skall åtala ?
det är här vi verkligen kommer i problem .
vems ansvar är det när det rör sig om ett organ som överskrider så många gränser ?
vi måste också ta hänsyn till medlemsstaternas oro .
förslaget att etablera en europeisk allmän åklagarmyndighet är mycket känsligt .
vi är alla medvetna om att en helhjärtad federalistisk inställning och en situation där en europeisk juridisk myndighet står över de nationella juridiska myndigheterna enligt vissa är att gå för långt .
men diskussionen måste starta och vi uppmanar därför regeringskonferensen att inleda diskussioner .
det viktigaste för parlamentet , i egenskap av europeiska unionens budgetövervakare , är hur man skall handskas med anställda inom europeiska unionens institutioner .
i en tid då vi ser över hela reformprocessen är det avgörande att vi ger rätt signaler .
människor måste inse att om de begår bedrägerier kommer de att åtalas , så är inte fallet för närvarande .
hela frågan om vi har laglig befogenhet att göra detta har palacio skisserat .
jag skulle vilja slå fast att min grupp kommer att föreslå en ändring som innebär att passusen om hur kommissionen bör handskas med denna fråga tas bort .
vi är medvetna om att detta är en känslig debatt .
vi vet att kommissionen kanske behöver spelrum för att förhandla fram en situation som alla parter kan acceptera .
låt mig bara göra klart att vi inte förbinder oss till en corpus juris här , inte förbinder oss till en europeisk allmän federal åklagare .
men vi förbinder oss definitivt att förändra ett status quo som är helt oacceptabelt .
herr talman ! jag skulle vilja börja med att lyckönska fru theato till hennes betänkande .
jag anser att det är ett utmärkt betänkande och att den övervägande delen av det kommer att stödjas av min grupp .
men jag får en stark känsla av att hon på detta stadium egentligen hade velat gå ett steg längre .
när jag lyssnat till diskussionerna under de senaste fem , sex månaderna skulle det mycket väl kunna vara fallet .
vi vet alla att vi 1995 kom överens om att man måste sörja för ett bättre straffrättsligt skydd för unionens ekonomiska intressen .
men medlemsstaterna var inte med på noterna .
det är helt enkelt ett politiskt faktum , och enligt vad jag tror kan vi för närvarande inte göra mycket åt detta .
den möjlighet som nu finns är att kommissionen på grundval av artikel 280 i fördraget tar nya initiativ , och jag skulle vilja föreslå kommissionen att verkligen göra detta så snabbt som möjligt .
min grupp är , i motsats till föregående talare som redan försvunnit , en stark förespråkare för en europeisk allmän åklagare .
min kollega jan-kees wiebenga kommer utan tvivel att ytterligare gå in på detta , för han har tidigare författat ett betänkande i ämnet .
det som vi har behov av , tror jag , är en definition på europeisk nivå av vad som exakt menas med bedrägeri och oegentlighet .
jag var själv med i undersökningskommittén om transittrafiken .
ett av de stora problemen på det området var att om man gör något fel , och då handlar det framför allt om europeiska unionens inkomster , så är det en oegentlighet i det ena landet och ett brott i det andra landet .
så kan vi inte ha det längre tyckte jag , i synnerhet inte för närvarande .
en allmän politisk punkt .
något som vi också kan konstatera i fråga om europavalet är att det låga valdeltagandet är ett faktum .
vi kan förbättra detta genom att snabbt ta itu med brottsligheten i europa , och det måste ske på europeisk nivå .
herr talman ! även mitt tack går till föredraganden .
theatos betänkande kan bidra till att det åter skapas förtroende för de europeiska institutionerna .
jag tror att vi alla verkligen behöver det , om vi tänker på resultaten från de senaste europavalen , och på valdeltagandet .
det är ju samma problem varje år .
revisionsrätten offentliggör sin rapport , och i rapporten beskylls medlemsstaterna för olika bedrägerier .
men de europeiska institutionerna har hittills haft alltför få möjligheter att ingripa och se till att något verkligen görs , att det avhjälps .
just detta förfarande minskar förtroendet varje år på nytt .
jag tror att theatos betänkande och hennes förslag kan bidra till att situationen vänder , och att det klargörs att de europeiska institutionerna ser till att de europeiska pengarna också satsas målinriktat och att det här inte förekommer några bedrägerier .
det är viktigt att vi efter det första steget som redan tagits , nämligen att ur uclaf skapa olaf , en oberoende institution , nu tar ett andra steg och även skapar en rättslig ram för olaf , så att olaf kan agera inom en säker rättslig ram .
till detta behöver vi den europeiska åklagarmyndigheten , som ser till att det finns en klar rättslig garanti , även för de misstänkta .
jag måste dock säga att min grupp tyvärr inte kommer att rösta enhälligt för ert betänkande .
jag hoppas att debatten kommer att övertyga ytterligare några personer .
betänkligheterna är tyvärr fortfarande alltför stora för att det här kommer att skapas en europeisk institution , som minskar subsidiariteten .
men jag vill bidra med min del så att theatos betänkande skall få ett större stöd .
herr talman ! vi är i allt väsentligt positiva till den resolution som lagts fram även om vi anser att detta inte kan bli annat än en uppmaning från parlamentet till rådet att genom en ändring av fördragen se till att skapa ett effektivt straffrättsligt skydd för unionens ekonomiska intressen .
inrättandet av en europeisk åklagare och tillskapandet av brottsrubriker som är gemensamma för samtliga länder inom unionen är utan tvekan en god idé , men jag anser det vara omöjligt att försöka förverkliga den utan att först ha inrättat en gemensam rättsordning för unionen .
vi talar ju här om straffrätten , det område där motståndet från nationalstaterna mot gemensamma regler är och alltid har varit starkt .
det är i själva verket otänkbart att man skulle kunna skapa gemensamma straffrättsliga regler för en enda sektor , nämligen skyddet av ekonomiska intressen , utan att först ha skapat ett gemensamt europeiskt rättssystem .
det räcker att man läser de exakta och uttömmande motiven i theatos betänkande för att man skall inse vilka problem som återstår att lösa .
men idén bör uppmuntras och det råder ingen tvekan om att man under dessa försök att skydda de ekonomiska intressena upptäcker behovet av att inrätta en gemensam corpus juris och att införa den i fördragen .
för egen del och som företrädare för min grupp vill jag också framföra en förhoppning om att unionens ekonomiska intressen blir en vägröjare för insikten om att det behövs ett europeiskt rättssystem som respekterar medborgarnas garanterade rättigheter , dvs. ett rättssystem som lyfter fram de garantier som , dessvärre , i många medlemsstater inte har nått upp till en godtagbar nivå .
jag uttrycker därför , som företrädare för min grupp , min uppskattning av theatos betänkande . men jag anser att det i grunden handlar om en fråga som måste föras upp på dagordningen för regeringskonferensen .
herr talman ! i betänkandet av theato om skyddet av europeiska unionens ekonomiska intressen föreslås bl.a. att man , i första hand , skall centralisera de straffrättsliga processerna genom att inrätta en europeisk åklagarmyndighet .
detta förslag står helt uppenbart i strid med andan i det nuvarande systemet , där straffrätten och straffrättsliga processer - centrala element i de nationella rättssystemen - skall lyda under varje folks suveränitet och varje stats exklusiva ansvarsområde .
idén om en europeisk åklagarmyndighet syftar tvärtom till att på sikt begränsa staterna och ge dem en underordnad roll i de här frågorna .
dessutom skulle förslaget utlösa en räcka reformer som är helt omöjlig att förutse .
enligt theatobetänkandet skulle en europeisk åklagarmyndighet vara nödvändig , bl.a. för att förbättra ledningen av undersökningarna vid byrån för bedrägeribekämpning , olaf .
men samtidigt får vi veta , i betänkandet av van hulten som diskuteras i dag , att den europeiska åklagarmyndigheten själv skall övervakas av en domstol i europeiska unionen .
på så sätt kan en liten europeisk reform dölja en medelstor , och en medelstor dölja en stor .
och då räknar jag inte med att en stor reform i sin tur kan dölja en gigantisk reform , eftersom vi snart kommer att få se ett förslag till en europeisk straffrätt och varför inte - på sikt - en europeisk justitieminister som kontrolleras genom en utvidgning av europaparlamentets befogenheter .
jag tror således att vi borde reflektera över den maktbalans som man riskerar att kullkasta genom att presentera reformer av det här slaget , vilka kan framstå som avgränsade .
slutligen anser vi att den här typen av förslag , såsom förslaget om en europeisk åklagarmyndighet , avslöjar en oförmåga att föreställa sig europa på något annat sätt än i en pyramidisk och centraliserad form , organiserad kring en överstat .
gruppen nationernas europa vill tvärtom ha ett europa med många centra som binder samman nationerna i ett nätverk .
detta nät skulle t.ex. kunna innebära en bättre samordning mellan nationella åklagarmyndigheter , och man skulle eventuellt kunna inrätta nationella utbildningar med inriktning på brott som skadar gemenskapens finanser . herr talman !
det finns således redan en juridisk struktur , och dess principer är bra .
vi behöver endast fullända den .
herr talman ! theato föreslår en institutionell revolution av två skäl .
allmänheten påstås vara likgiltig inför 20 miljoner arbetslösa och tusentals galna kor , men oroad över de bedrägerier som äventyrar de ekonomiska intressena , och dessa två skäl skulle motivera två bestämmelser : en europeisk straffrätt om anti-gemenskapliga förbrytelser och en europeisk allmän åklagarmyndighet .
theato har förresten , sannolikt , glömt ett europeiskt fängelse , eftersom fbi - den europeiska polisen - existerar i och med olaf .
allt detta skulle inrättas genom två förordningar , en för åklagarmyndigheten och en för straffrätten .
det är förordningar som antas på grundval av artikel 280 i fördraget , dvs. med utgångspunkt i den avledda rätten , för det som utmärker den avledda rätten är att man tillåter alla strömningar som leder i andra banor .
det finns faktiskt två strömningar .
först och främst den klassiska ideologiska , eurofederalistiska strömningen : för en gemensam marknad , en gemensam mervärdesskattesats , en gemensam diplomati , en gemensam armé och nu en gemensam straffrätt och en gemensam åklagare .
allt detta för att bekämpa bedrägerier som underskrider en miljard euro , samtidigt som man mister tiotals miljarder euro på grund av allmänna preferenssystemet , frihandelsområdena , tullgåvor till chiquita och miljarder som förlorats på den fjärde resursen , bni , ett resultat av pakten om finansiell åtstramning .
sedan har vi den puritanska strömningen ; det nordtyska europa , det lutheranska och calvinistiska europa , kväkareuropa , som vill påtvinga oss sin moraliska ordning .
för i grunden är det så , att ju mer man lättar på seder och bruk , desto hårdare håller man i plånboken .
herr talman , mina damer och herrar ! det är absolut nödvändigt med ett verksamt straffrättsligt skydd för europeiska unionens intressen , i dag mer än någonsin .
bedrägeri- och korruptionsskandalerna i det förflutna har på lång sikt skakat förtroendet hos europas medborgare .
trovärdigheten i de ansträngningar vi gör här i parlamentet för att de ekonomiska medlen skall satsas korrekt står och faller med våra ansträngningar för att behandla dem och förhindra dem i framtiden .
hit hör inte bara administrativa , utan också strukturella förändringar , dvs. vi måste skapa de instrument med vilka man över huvud taget kan garantera ett straffrättsligt skydd .
regeringskonferensen 2000 är lämplig som diskussionsforum för detta .
nu kan man naturligtvis inta den ståndpunkten att straff- och straffprocessrätten hör till medlemsstaternas rättssystem och inte kan röras när man har en subsidiaritetsprincip .
själv hör jag utan tvivel till dem som förfäktar denna princip och till motståndarna av all vidare utvidgning av de europeiska ansvarsområdena .
just i samband med kraven på regeringskonferensens arbete bör tyngdpunkten ligga på att fordra en klar ansvarsavgränsning .
men detta innebär inte någon motsägelse , ty när man kräver ett straff- och straffprocessrättsligt instrument , så som anförs i betänkandets rekommendation i och ii , handlar det egentligen om att iaktta eu : s ursprungliga egna intressen , som såtillvida inte skadar medlemsstaternas rättsliga intressen , utan tvärtom stöder dem , åtminstone indirekt .
förenligheten med de olika nationella rättssystemen , som bekräftats av experterna , visar att man i europa har mycket gemensamt även på det straffrättsliga området , exempelvis när det handlar om innehållet i de här tillämpliga åtalspunkterna .
med hänsyn till dessa synpunkter anser jag att skapandet av en sådan ram som krävts är riktigt och också är påbjudet som en vidareutveckling av olaf .
herr talman ! kommer en europeisk offentlig åklagare att kunna avskaffa fotbollsbedrägerierna med eu-medel ?
vi kan istället komma långt med de befintliga instrumenten .
eurojust skulle kunna vara ett alternativ till den europeiska offentliga åklagaren , vilket föreslogs på det senaste toppmötet .
eurojust skall i inledningsskedet lyda under europol och stödja forskningen i brottsfrågor .
det är precis ett sådant praktiskt samarbete det finns behov av .
olaf , europol och konventionen om utlämning och ömsesidig rättshjälp skall utnyttjas fullt ut , och när bedrägerikonventionen från 1995 slutligen blir ratificerad av medlemsstaterna , kan vi även komma långt med hjälp av den .
jag håller emellertid med föredraganden : det är fullständigt oacceptabelt att de flesta medlemsstaterna ännu inte har ratificerat den .
det är helt enkelt för dåligt och jag förstår mycket väl att folk blir otåliga och kräver att vi i stället skall få en gemensam europeisk åklagare .
det är emellertid en stor mastodont att bygga upp .
det är ändå bara de grövsta fallen som kommer att få straffrättsliga konsekvenser .
90 procent av fallen kommer att utgöra disciplinfrågor om försummelse eller inkompetens .
i stället finns det behov av en ordentlig intern kontroll och bättre möjligheter att avskeda folk .
vi skall ändra tjänsteföreskrifterna och det disciplinära förfarandet och inte minst skall vi ändra praxis .
för närvarande används aldrig artikel 52 i tjänsteföreskrifterna om avskedande på grund av grov försummelse .
skall vi inte se till att rensa upp ordentligt och hålla rent framför vår egen dörr , innan vi förhastar oss och börjar bygga upp nya förkromade institutioner ?
herr talman ! vi vill allesammans gärna göra något för den europeiska bedrägeribekämpningen .
men frågan är nu : gör europeiska unionen också något för denna ?
svaret är att vi vet alldeles för litet om detta .
toppmötet i tammerfors handlade om brottsbekämpning .
alla var så kallat nöjda med detta , men i själva verket gjordes det inte några större framsteg .
det finns fortfarande ingen gällande europeisk antibedrägerilagstiftning , eftersom medlemsstaterna , vilket redan har sagts , inte har ratificerat de framlagda fördragstexterna .
på det området måste det således hända mycket .
och vad är det då som måste hända ?
det är två saker , och i theatos betänkande framkommer detta på ett klart och tydligt sätt .
för det första , i alla europeiska unionens medlemsstater måste samma straffbestämmelser gälla i fråga om europeiskt bedrägeri .
likriktning på detta begränsade område .
för det andra måste verkligen en europeisk åklagarmyndighet inrättas , och den skall ha två uppgifter : för det första att stödja de nationella allmänna åklagarna , att hjälpa till med åtal i fråga om europeiska bedrägerimål , och för det andra att övervaka europol och olaf i rättsligt avseende , för detta är två utredande myndigheter som för närvarande kan operera okontrollerat i rättsligt avseende .
den europeiska åklagarmyndigheten är inte någonting att vara rädd för ; det jag hör här runt omkring mig är bara skräckscenarior .
det är helt enkelt något mycket positivt , precis som europol .
europol , polissamarbetet , står inte över de nationella polismyndigheterna , utan finns med tanke på informationsutbytet mellan polismyndigheterna .
det är precis på det sättet som en liten begränsad europeisk åklagarmyndighet måste börja arbeta . det gäller inte bara under uppspårningsfasen , utan också under åtalsfasen .
parlamentet är för detta .
den oberoende expertkommittén är för detta .
jag uppmanar ministerrådet och europeiska kommissionen att också erkänna denna åtgärd .
herr talman ! jag skall koncentrera mig på frågan om corpus juris .
jag vill verkligen stödja det morgan sade om detta .
corpus juris är någonting som sattes ihop utan någon offentlig debatt eller deltagande alls .
tanken med en europeisk allmän åklagare med överordnad jurisdiktion inom eu : s territorium skulle få stora konsekvenser för de traditionella systemen både i irland och i storbritannien .
planerna på en enda strafflagstiftning och en europeisk allmän åklagare är någonting medlemsstaterna har rätt att få information om .
när planen först gjordes upp sade de att den skulle vara begränsad till fall av bedrägeri mot eu : s budget .
men när corpus juris lanserades i san sebastian 1977 - inför en mycket utvald publik på 140 jurister , utan inbjudna media - sade den dåvarande talmannen i europaparlamentet , gil-robles gil-delgado , att han ansåg att den var på embryostadiet och att avsikten var att utvidga eu : s befogenheter på brottsmålssidan till att omfatta all kriminell verksamhet .
vi behöver en offentlig debatt om detta .
medlemsstaterna och medborgarna i medlemsstaterna måste få ordentlig information .
frågan om hotet mot det traditionella juridiska systemet i irland och storbritannien måste tas upp .
det behövs mycket större öppenhet och insyn än hittills i denna fråga .
det är oacceptabelt att någonting dylikt har prackats på eu : s medlemsstater utan någon ordentlig offentlig debatt .
herr talman , kära kolleger ! i budgetkontrollutskottet avstod jag från att rösta om denna text i min egenskap av företrädare för de radikala ledamöterna , för jag delar den oro som på ett så kunnigt vis formulerats av företrädaren för en annan mycket viktig juridisk tradition , dvs. den som har formen av common law .
med den här texten rör vi oss verkligen i utkanten av vad som är möjligt , eftersom vi anser att det finns frågor som måste lösas och att det är viktigt att bedrägerierna inom gemenskapen stoppas , att de stryps .
men det sätt på vilket vårt utskott , tack vare ordföranden theatos energi och envishet , har för avsikt att förverkliga intentionerna i denna text får inte ske utan kritik .
en annan viktig kritik som kan riktas mot texten gäller sekundärrätten .
artikel 280 i fördraget ger rådet rätt att bestämma om lämpliga instrument för att bekämpa bedrägeriet .
men vi blir ändå en aning förvånade över att man vill inrätta en institution , vilket innebär ett kvalitetssprång , utan att genast kunna förutse vilka motåtgärder som kommer , dvs. man bortser från försvaret och därmed möjligheten att åklagare och försvarare skall kunna fungera effektivt i ett så viktigt rättssystem .
genom att avstå från att rösta i utskottet har vi velat uttrycka denna vår tveksamhet .
herr talman ! jag tror att det är något som måste sägas tydligt i denna fråga i denna församling , i plenarsammanträde och i utskotten , eftersom det är uppenbart att debatten inte får bortse från den kulturella bakgrunden , den juridiska kulturen och de miljöer i vilka de institutionella frågorna skall tas upp .
vi står inför mycket allvarliga händelser som i det förflutna verkade vara en tradition .
i dag har något förändrats , åtminstone när det gäller mekanismerna , framför allt när det gäller kontrollen , men vi är ändå inte nöjda , framför allt inte om man i berörda fora pratar om en europeisk åklagare , brott , bedrägerier , förskingring och avslöjanden av hemligheter på europeisk nivå .
jag anser naturligtvis att vi måste skydda gemenskapens intressen och dess rykte , förutom relationerna med bidragsgivarna , som utgör en omistlig och avgörande del av gemenskapens liv .
av den anledningen är det riktigt att undersöka frågan om ett skydd av intressen av mer allmän och universell natur , och att på ett bättre sätt förena sig med rättssystemen inom de enskilda staterna .
i det sammanhanget uppstår en känsligare fråga : hur förhåller sig en europeisk åklagare till de enskilda medlemsstaterna och det rättssystem som är uppbyggt inom ramen för dem ?
detta är en fråga som fortfarande måste tas upp såväl ur kulturell som praktisk synpunkt .
i dag riskerar vi att lägga en ny institution ovanpå de många skilda institutioner som redan existerar i de enskilda länderna .
herr talman ! jag vill gärna helt snabbt säga något om två punkter .
för det första : jag vill inte referera till de filosofiska frågorna om medlemsstaternas subsidiaritet och suveränitet , även om jag absolut anser att en sådan debatt bör föras , eftersom mitt regelbundna tittande på brittiska tv-sändare ändå får mig att inse vad nationella politiker där betraktar som ett hot mot den inhemska rättskulturen från kontinentens sida .
ibland är det nästan kabarébetonat och förtjänar att diskuteras . men det är inte det jag vill tala om .
jag vill tala om theatos betänkande .
jag tror att man har trasslat in sig i de juridiska svårigheter som finns här - och uppenbarligen finns det bara en mycket liten möjlighet för europeiska unionen att ta upp dessa åtalspunkter som europeiska åtalspunkter .
jag refererar till rekommendationerna 1 och 2 .
det står ju där inte längre något om en europeisk åklagare , utan av juridiska orsaker har det nu blivit en oberoende europeisk myndighet , med theatos ord tidigare en organism .
där har vi uppenbarligen problem med den rättsliga grunden .
sedan har vi problem med åtalspunkterna .
det har inte ändrats .
där finns det fortfarande åtalspunkter , som så att säga också går utöver de europeiska åtalspunkterna , eller åtminstone kan gå utöver dem , exempelvis penningtvätt , häleri och stämpling .
i det avseendet anser jag att det finns juridiska oklarheter , som bör undanröjas .
men det som är absolut nödvändigt , och därför kommer vi att rösta för punkt 1 utan dessa rekommendationer , är en klar politisk signal från parlamentet till kommissionen och rådet att vi med hjälp av en klar rättsakt vill ha ett slut på de förhållanden , som har gripit omkring sig .
herr talman ! parlamentet har sedan flera år krävt en specifik och enhetlig straffrätt till skydd för unionens ekonomiska intressen .
sanningen är att frustrationen ökar när vi konstaterar svagheterna i konventionen ( och protokollen i anslutning till detta skydd ) , som fem år efter att den undertecknats ännu inte har ratificerats eller trätt i kraft .
mer voluntaristiska försök , som det nuvarande olaf , övervinner inte den legitima oron över garantisystemet för de individuella rättigheterna .
förslagen i theatos betänkande för att uppmuntra kommissionen att lägga fram en rättsakt om straffrättsliga bestämmelser till skydd för unionens ekonomiska intressen med typfall för brott , framför allt oredlighet avseende bidrag från och avgift till gemenskapens budget , är enligt vår mening ett försök att införa en ny och allt nödvändigare enhetlig straffrätt i gemenskapen .
samtidigt är de en vädjan om inrättande av ett &quot; oberoende europeiskt organ &quot; , som samordnar och kontrollerar att olaf : s utredningsverksamhet följer gällande bestämmelser , utan att det påverkar medlemsstaternas rättskipning och under eg-domstolens övervakning .
slutligen , i tammerforsbeslutens fotspår tas i betänkandet återigen ett europeisk åklagarämbete upp , vilket kommissionär antónio vitorino i ett lämpligt ögonblick beslutade sätta ljuset på genom att begära att regeringskonferensen skulle ta upp skapandet av denna nya tjänst i sin dagordning , det ämbete som alla i dag anser är nödvändigt .
eftersom behovet av rättslig och effektiv disciplin i institutionerna vidhålls , genom att tillsluta unionens ekonomiska system med en europeisk materiell och processuell rätt anpassad till förtroendet för gemenskapens ekonomiska liv , stöder vi detta betänkande .
emellertid finns det några mycket enkla frågetecken .
finns det tillräckligt med rättslig grund för att motivera skapandet av en ny specifik straffrätt för gemenskapen som , även om man kan kalla den subsidiär , i praktiken och i vissa områden alltid kommer att strida mot medlemsstaternas traditionella och partiella straffrätt ?
skulle det inte vara mer politiskt korrekt , när det råder tvivel , att föra upp reformen av rättssystemet på regeringskonferensens dagordning , och alltså ta upp dessa förslag i den mer allmänna reformen av unionens rättssystem , och ta upp dem i den bild man vill ge den europeiska åklagaren ?
är inte dessa frågor av största intresse för en revidering av fördragen som kan bidra till att befästa området med frihet , säkerhet och rättvisa i unionen ?
herr talman ! eu utsätts i dag för hård granskning .
förtroendet för unionen är allvarligt skadat .
för att råda bot på detta krävs krafttag .
vi välkomnar därför ökade resurser till olfaf , så att vi effektivare kan utreda alla misstankar .
vi ser det samtidigt som självklart att de som begår brott mot eu på ett effektivt sätt måste kunna ställas till ansvar .
det är beklagligt att konventionen om skydd för unionens ekonomiska intressen har genomförts i så få medlemsstater .
vi menar därför att det är rimligt att kommissionen får i uppdrag att lägga fram förslag , som innebär att den rättsliga ram som redan finns vidareutvecklas .
däremot är jag inte övertygad om att en sådan effektivisering kräver en gemensam europeisk lagstiftning eller en centralisering av sådan brottsbekämpning .
i dagsläget är jag därför skeptisk till idén om en europeisk åklagare , vilken knappast är möjlig att genomföra inom ramen för dagens fördrag .
vi tror mer på eurojust , där nationella åklagare samarbetar .
det stora problemet är inte att brott mot unionen inte beivras , utan att de så ofta begås och alltför sällan upptäcks .
utmaningen för kommissionen och för oss är dock att finna rätt mix .
de bedrägerier och den misshushållning som förekommer får inte leda till att vi fastnar i en ålderdomlig hierarkisk byråkrati , som genom överdriven detaljkontroll förhindrar utvecklingen av modern förvaltning .
därför välkomnar vi den offensiva synen i van hultenbetänkandet .
huvudlinjen bör vara att varje förvaltning tar ansvar för sin egen kontroll .
våra erfarenheter av modern förvaltning säger oss att öppenhet , decentralisering av ansvaret och kvalificerad utvärdering ofta är lika effektivt som byråkratisk detaljkontroll .
den stora utmaningen är därför att skapa en modern och effektiv förvaltning utan att förlora i rättssäkerhet och kontroll .
det kräver personalutbildning , modernare rekryteringsmetoder och framför allt öppenhet och insyn .
att kunna granska förvaltningen effektivt är det bästa skyddet mot oegentligheter .
tack , kommissionär schreyer .
heaton-harris ( ppe-de ) .
( en ) herr talman ! som en ordningsfråga skulle jag vilja be er om ett klargörande av arbetsordningen , nämligen artiklarna 133.2 och 138.4 .
de handlar båda om omröstning .
är det inte så att vid andra omröstningar än omröstningar med namnupprop skall omröstning först ske genom handuppräckning och först sedan , om det finns tvivel om utgången , skall vi använda det elektroniska voteringssystemet ?
det stämmer att jag genomförde en omröstning med handuppräckning , eftersom ingen grupp hade begärt en omröstning med namnupprop .
som ni vet genomförs endast omröstningar med namnupprop och elektroniska omröstningar om kollegerna begär detta .
i det här fallet kan jag försäkra er att det fanns en överväldigande majoritet för det direktiv som vi just har röstat igenom .
herr talman , jag syftade inte på just denna omröstning utan på omröstningar i allmänhet .
det är uppenbart att vissa ordförande inte tittar på händerna , så att säga , utan går direkt till det elektroniska voteringssystemet .
jag undrade om detta är ett korrekt tillvägagångssätt .
jag vet att det tar längre tid , men borde vi inte alltid först räcka upp händerna ?
jag försäkrar er , kära kollega , att jag kommer att vara mycket uppmärksam på hur många händer som räcks upp .
jag hoppas att det blir många då det är dags för omröstning .
förslag till europaparlamentets och rådets direktiv om tillnärmning av medlemsstaternas lagstiftning om märkning och presentation av livsmedel samt reklam för livsmedel ( kodifierad version ) ( kom ( 1999 ) 0113 - c4-0212 / 1999 - 1999 / 0090 ( cod ) ) ( utskottet för rättsliga frågor och den inre marknaden )
förslag till rådets förordning ( eg , euratom ) om genomförande av beslut 94 / 728 / eg , euratom om systemet för gemenskapernas egna medel ( kodifierad version ) ( kom ( 1997 ) 0652 - c4-0018 / 98 - 1997 / 0352 ( cns ) ) ( utskottet för rättsliga frågor och den inre marknaden )
betänkande ( a5-0106 / 1999 ) av varela suanzes-carpegna för fiskeriutskottet om förslag till rådets förordning om slutande av det protokoll i vilket de fiskemöjligheter och finansiella motpartsmedel fastställs som föreskrivs i avtalet mellan europeiska ekonomiska gemenskapen och demokratiska republiken são tomé och príncipes regering om fiske utanför são tomé perioden 1 juni 1999 - 31 maj 2002 ( kom ( 1999 ) 0550 - c5-0305 / 1999 - 1999 / 0228 ( cns ) )
andrabehandlingsrekommendation ( a5-0105 / 1999 ) från utskottet för regionalpolitik , transport och turism om rådets gemensamma ståndpunkt inför antagandet av europaparlamentets och rådets direktiv om harmonisering av examineringskraven för säkerhetsrådgivare för transport av farligt gods på väg , järnväg eller inre vattenvägar ( c5-0208 / 1999 - 1998 / 0106 ( cod ) ) ( föredragande : koch )
det är med stor tillfredsställelse jag välkomnar detta betänkande om en bättre harmonisering inom utbildningen av säkerhetsrådgivare för transport av farligt gods .
under de senaste åren har de nationella och internationella transporterna av farligt gods ökat avsevärt , vilket har ökat olycksriskerna .
vissa av olyckorna har berott på en otillräcklig kunskap om de risker som hänger samman med den här typen av transporter .
det har således visat sig nödvändigt att anta åtgärder - inom ramen för genomförandet av den inre marknaden - för att ombesörja ett bättre förebyggande av risker .
genom direktiv 96 / 35 / eg uppfylldes det kravet .
följaktligen har de företag som transporterar farligt gods och de företag som genomför lastning och lossning i samband med sådana transporter med rätta sett sig tvingade att respektera regler om riskförebyggande , vare sig det gäller transporter på väg , järnväg eller inre vattenvägar .
för att göra det lättare att förverkliga detta mål , föreskrev direktiv 96 / 35 / eg att de säkerhetsrådgivare som utses för transporter av farligt gods skall ha en lämplig yrkesutbildning .
målet med denna yrkesutbildning för rådgivare skulle vara en kunskap om de viktigaste lagar , förordningar och bestämmelser som gäller för dessa transporter .
detta utgjorde ett framsteg för några år sedan , men så småningom uppstod problem eftersom det saknas specifika bestämmelser om harmoniseringen av examineringsvillkoren .
det föreföll därför nödvändigt att komma tillrätta med den svagheten , för att nå en högre och enhetlig utbildningsnivå för säkerhetsrådgivare , men också för att undvika skillnader mellan utbildningskostnader och följaktligen en inverkan på konkurrensen mellan medlemsstaternas företag .
kommissionens förslag syftar till att garantera en enhetlig utbildning av säkerhetsrådgivarna .
förslaget avgränsar minimiinnehållet i en examen och fastställer den behöriga myndighetens uppgifter , såväl som vilka krav som skall uppfyllas av examineringsorganen .
parlamentet har ställt sig positivt till denna text .
men det har ändå lagt fram flera ändringsförslag , varav de flesta har införlivats i rådets gemensamma ståndpunkt , t.ex. att det skall vara nödvändigt att genomföra en fallstudie och ge utlåtande om tillstånd till vissa dokument inom ramen för en &quot; specificering av de examineringsformer som examineringsorganet föreslår &quot; .
jag ger för övrigt mitt stöd till att tidsfristen för genomförandet av dessa bestämmelser skjuts upp till tre månader efter det att direktivet har trätt i kraft , med hänsyn till vad som är realistiskt .
jag vill avsluta genom att insistera på det faktum att rådgivarnas yrkeskvalifikationer kommer att bidra till en förbättrad servicekvalitet till användarnas fördel , och det kommer att minimera de olycksrisker som en försämrad miljö kan medföra liksom de allvarliga skador vilka kan skada den fysiska integriteten hos alla de personer som kan komma i kontakt med farligt gods .
betänkande ( a5-0104 / 1999 ) av koch
i oktober förra året uttalade jag mig om hatzidakisbetänkandet om transport av farligt gods på järnväg .
mina synpunkter i dag står inte långt ifrån dem jag hade då .
de kan sammanfattas på följande sätt : jag beklagar att vi ständigt skjuter upp antagandet av harmoniserade normer på ett så avgörande område som transport av farligt gods . det skadar människors säkerhet och miljön .
jag vill erinra om att ett direktiv om tillnärmning av medlemsstaternas lagstiftning om transport av farligt gods på väg trädde i kraft den 1 januari 1997 .
det innehåller ett antal övergångsbestämmelser som var giltiga fram till den 1 januari 1999 .
från och med det datumet borde vi ha uttalat oss om ett förslag från europeiska kommissionen , med syftet att få dessa undantag att upphöra .
enligt det nuvarande förfarandet är det europeiska standardiseringskommittén ( cen ) som föreslår normer på det här området . dessa upptas sedan i europeiska överenskommelsen om internationell transport av farligt gods på väg , som undertecknades i genève 1957 ( mer känt under förkortningen adr ) och tillämpas i hela europa , och vars bestämmelser utgör grunden för den lagstiftning som är tillämplig i europeiska unionen .
men cen har inte kunnat utföra sitt arbete inom den anvisade tiden .
syftet med det förslag från kommissionen som vi diskuterar i dag är därför att ändra på direktivet för att lösa problemen på kort sikt , och inte att sätta punkt för övergångssystemet , vilket borde ha varit fallet !
precis samma sak hände när det gällde transport av farligt gods på järnväg , fast med en skillnad : en tidsfrist fastställdes .
i dag har vi inte den blekaste aning om när cen kommer att kunna ge oss konkreta förslag .
fram till dess är det egentligen onödigt för medlemsstaterna att ändra sina nationella bestämmelser .
i betänkandet accepteras också att man inför en viss flexibilitet , och man tillerkänner staterna möjligheten att anta eller tillämpa olika normer .
medlemsstaterna skulle således kunna fortsätta att tillämpa sina egna normer för vissa transportabla tryckbärande anordningar , eftersom de europeiska normerna inte är tillräckliga i det fallet .
staterna kan också anta olika bestämmelser för transporter av lokal art och enstaka transporter .
med denna röstförklaring vill jag i dag uttrycka mitt djupa missnöje och min stora oro .
betänkande ( a5-0108 / 1999 ) av schroedter
herr talman ! jag skulle vilja lägga tyngd bakom min röstförklaring genom denna muntliga förklaring med anledning av schroedterbetänkandet om den regionala utvecklingen .
jag vill uppmana såväl medlemsstaterna som kommissionen att ägna tillräcklig uppmärksamhet åt de stora välfärdsskillnader som finns kvar mellan de olika regionerna i europa .
det gäller inte bara skillnaden i inkomst per capita , utan det är framför allt de stora skillnaderna beträffande sysselsättning som fortsätter att vara en källa till oro .
trots det faktum att gemenskapen , bland annat via strukturfonderna , lägger ned avsevärda summor på att bekämpa skillnaderna mellan chanserna till utveckling för våra regioner i europa kvarstår dessa skillnader .
det gör att jag ställer mig frågan om inte gemenskapen bör lägga om kursen på ett mer drastiskt sätt , och på grundval av mycket strikta utvärderingar bör övergå till en kursändring och till en ändring av målsättningarna som gör det möjligt att bedriva en effektivare kamp mot skillnaderna i välfärd och sysselsättning .
herr talman ! vad gäller schroedters betänkande är jag medveten om , och har fått bekräftat av barnier , att reglerna om komplementaritet vad strukturfonderna beträffar bara kan tillämpas på medlemsstatsnivå och inte är tillämpliga på ett transitivt och öppet sätt inom medlemsstaterna till förmån för självstyrande regioner såsom wales eller skottland .
jag tycker att detta är mycket otillfredsställande .
jag hoppas att vi kan ompröva denna fråga vid ett senare tillfälle .
jag vill göra klart att jag har denna viktiga invändning även om jag röstade för betänkandet .
. ( en ) i schroedters betänkande talar man om behovet att främja partnerskap vad beträffar ianspråktagandet av eu : s strukturfonder för perioden 2000-2006 .
jag anser att detta är särskilt viktigt eftersom medlen i eu : s strukturfonder alltid används på ett sätt som maximerar olika regioners ekonomiska utveckling när lokala och regionala myndigheter är involverade i beslutsfattandet om hur dessa fonder skall användas .
i egenskap av ledamot av europaparlamentet för leinsters valkrets har jag alltid hävdat behovet av att förverkliga lokala initiativ som stöds av nationella eu-fonder .
jag anser att den irländska regeringen och europeiska kommissionen och olika eu-regeringar inte själva kan besluta om specifika utgiftsprioriteringar .
jag anser att lokala myndigheter och grupper från den privata sektorn och frivilligsektorn bör vara fullt involverade i beslutsfattandet om hur de europeiska strukturfonderna skall användas .
vi har till exempel sett vilken framgång programmen leader i och ii har haft i irland i form av de arbeten som har skapats genom dessa program på den irländska landsbygden och inom europa .
programmet leader iii skall verkställas någon gång senare i år .
kärnan i leader-programmet är att ge offentliga , privata och ideella grupper möjlighet att slå ihop sina resurser så att en permanent och hållbar sysselsättning skapas i små och medelstora företag på landsbygden .
detta är ett klassiskt exempel på hur partnerskapskonceptet fungerar , och sådana program måste ingå i dess befogenheter .
den europeiska fonden för fred och försoning har också varit framgångsrik när det gäller att skapa arbetstillfällen i irlands gränsområden .
även här finns ett aktivt deltagande från offentliga , privata och ideella grupper vilka lämnar förslag om hur särskilda fondmedel bäst kan användas för att understödja olika lokala projekt för att skapa sysselsättning i denna region .
under nästa runda för eu : s strukturfonder 2000-2006 kommer andra eu-initiativ såsom &quot; equal &quot; och &quot; urban &quot; att vara i full gång .
dessa initiativ måste också involvera för att identifiera var de europeiska strukturfonderna kommer bäst till nytta .
föredraganden hänvisar till behovet att skapa en samordnad inställning till planer och program för nya eu-strukturfonder .
de måste främja ett decentraliserat , effektivt och mångsidigt partnerskap grundat på kunskaperna och engagemanget inom regionala och lokala myndigheters alla sektorer .
detta är mycket känsligt eftersom avgörande ekonomiska och sociala problem i vårt land inte kan lösas om det inte finns en samordning av nationell , europeisk och lokal bidragsgivning .
detta betänkande föranleder följande fråga : vilket är regionalpolitikens existensberättigande ?
för att minska de regionala skillnaderna givetvis .
men det hänger framför allt samman med den europeiska marknaden , som a priori skall garantera oss en bättre fungerande ekonomi , men som också kan vara en källa till orättvisor .
jacques delors brukade säga att marknaden är närsynt , därav den politiska nödvändigheten av att minska skillnader .
det handlar om den solidaritet som är ursprunget till den europeiska sociala modell som vi alla försvarar , och som har gett upphov till den ekonomiska och sociala sammanhållningen .
det verkliga politiska målet , på samma sätt som när det gäller ekonomi och valutafrågor , är något som utvecklas i samarbete med medlemsstaterna , regionerna och de lokala myndigheterna . kommissionens uppgift är att med hjälp av riktlinjer visa medlemsstaterna vilken linje som skall följas , för att de eftersträvade målen skall uppnås inom ramen för programplaneringen .
därför kommer jag att stödja detta betänkande , samtidigt som jag beklagar , av skäl som har att göra med tidsplanen , att europaparlamentet inte rådfrågades förrän mycket sent i fråga om de riktlinjer som skall hjälpa medlemsstaterna , regionerna och de lokala myndigheterna med programplaneringen av mål 1 , 2 och 3 .
i övrigt önskar jag att kammaren också tar hänsyn till yttrandet från utskottet för sysselsättning och sociala frågor , vilket tillfogar en reflektionsplan för centrala frågor såsom bekämpningen av social utslagning , stödet till den sociala ekonomin och genomförandet av sysselsättningsstrategin .
schroedters arbete är ett steg mot en större öppenhet och effektivitet inom ramen för de strukturella stöden .
hon sätter värde på den växande och ytterst viktiga roll som samtliga aktörer har , och särskilt våra lokala partner - de enda som kan definiera specifika frågor och sociala problem .
därför vill vi försäkra oss om att de partnerskap som skall genomföras blir verkliga partnerskap , decentraliserade partnerskap som involverar samtliga berörda aktörer , och därför omformulerar vi vårt krav på att det skall inrättas ett centrum för förvaltning av strukturstöden i medlemsstaterna , med uppdraget att samordna genomförandet och förvaltningen av stöden .
för det ändamålet krävs det att utvärderingskommittéerna står öppna för europaparlamentets ledamöter , föreningar , näringsidkare som berörs av projekten samt det civila samhället .
dessa riktlinjer är ett steg för att göra gemenskapens strukturstöd effektivare .
ändras de enligt schroedterbetänkandet , går de i rätt riktning .
de uppmanar också till en allmän debatt om sammanhållningspolitikens framtid efter år 2006 , men det är en annan debatt .
låt oss stödja detta första steg i väntan på den .
. ( en ) i detta betänkande krävs drastiska nedskärningar av det illegala statliga stöd vissa medlemsstater delar ut .
även om jag helhjärtat stöder detta syfte skulle jag mycket hellre se att ett sådant stöd avskaffades helt .
enligt min mening är illegalt statligt stöd inte mycket bättre än statligt sponsrad social dumpning .
vi är alla emot social dumpning när förövaren är den välmående bilindustrin , då måste vi också vara emot den när förövaren är en regering .
om vi skall kunna få en effektiv inre marknad som gör den europeiska industrin konkurrenskraftig globalt och skapar välstånd och sysselsättning för alla européer måste vi ha en jämn spelplan .
illegalt statligt stöd däremot förstör konkurrenskraftiga företag och skapar arbetslöshet .
det finns förstås fall där statligt stöd kan vara nödvändigt och legitimt , för att till exempel hjälpa företag vid omstruktureringar .
i alla sådana fall måste dock strikta kriterier uppfyllas och tillstånd från europeiska kommissionen inhämtas i förväg .
oavsett om vi talar om nötkött till frankrike eller mutor till industrin får inte eu : s medlemsstater tillåtas att driva gäck med lagen .
jag stöder med entusiasm förslaget i betänkandet att offentliggöra en &quot; resultattavla &quot; som visar det statliga stödet per medlemsstat .
länder som hävdar att de ligger i europas hjärta men som systematiskt bryter mot dess regler bör demaskeras och deras hyckleri avslöjas .
medlemsstaterna kan inte tillåtas proklamera europeisk solidaritet offentligt och samtidigt försöka underminera den inre marknaden privat .
jag blir något uppmuntrad av det faktum att nivån på det statliga stödet till industrin i europa tycks minska .
emellertid återstår mycket att göra , och jag uppmanar kommissionen att vara mycket tuffare när den exponerar europas bidragsnarkomaner .
- ( pt ) eftersom kommissionens viktigaste instrument för att övervinna de regionala skillnaderna är strukturfonderna och sammanhållningsfonden , är det väsentligt att europaparlamentet deltar i utformandet av dess allmänna vägledande riktlinjer utan att det sker på bekostnad av subsidiariteten , då fastställande av utvecklingsstrategierna i varje land är medlemsstaternas sak .
tyvärr har europeiska kommissionen redan gått framåt med sina riktlinjer och parlamentets ståndpunkt är inte mycket värd för programmen under perioden 2000-2006 .
det är dock viktigt att trycka på betydelsen av att dessa fonder först och främst prioriterar utvecklingen i de länder och regioner som har störst svårigheter och i gemenskapens yttersta randområden , vilket portugal och regionerna azorerna och madeira är exempel på , för att uppnå ekonomisk och social sammanhållning .
i själva verket uppfyller inte kommissionens riktlinjer dessa mål helt .
det är också viktigt att det finns precisa indikationer och tillräckliga medel för att skapa kvalitativ sysselsättning med rättigheter liksom för att effektivt främja lika rättigheter och möjligheter , stödja en social och solidarisk ekonomi , landsbygdens utveckling , de små och medelstora företagarna , samt för att förbättra livskvaliteten för stadsbefolkningen i fattigare områden , främst inom området för bostäder som subventioneras med allmänna medel , för att härigenom uppnå en hållbar utveckling i städerna .
( it ) om innehållet i artikel 158 i eg-fördraget syftar till att främja en harmonisk utveckling av hela gemenskapen , så måste vi tyvärr konstatera att vi fortfarande är långt från målet att utjämna skillnaderna . det är till och med så , till exempel för de italienska områden som återförts till mål 1 , att skillnaderna paradoxalt nog ökar , framför allt på grund av att de lokala organisationernas förmåga att hantera gemenskapens rutiner fortfarande är bristfällig och att det råder ett permanent kaos när det gäller förvaltningen .
trots ingreppen i regelsystemet har vi ännu inte lyckats få gemenskapens strukturer att arbeta snabbare . om man inte förenklar byråkratin så blir det svårt att uppnå gemenskapens mål , som är att genomföra reformer präglade av effektivitet och koncentration .
i det avseendet är kommissionens dokument bristfälligt , eftersom här inte finns några som helst rekommendationer till medlemsstaterna om hur man skall kunna förenkla nationella regler och rutiner när det gäller hur de nationella myndigheterna skall presentera och informera om olika projekt , eller när det gäller finansiering , genomförande och kontroll .
små och medelstora företag , mikroföretag och hantverkare är fortfarande &quot; svaga subjekt &quot; , eftersom de hinder som finns i regler och byråkratiska rutiner i vissa medlemsstater , bland annat italien , just för dem gör det betydligt svårare att få tillgång till strukturfonderna .
ett viktigt handicap är regionernas och andras oförmågan och bristande möjligheter att planera i god tid , varför kommissionen , som på grundval av beslutet om riktlinjer 97 / 99 ( howittsbetänkandet ) hade kunnat rådfråga parlamentet i god tid , i själva verket hittade ett bekvämt alibi när man inrättade den förkortade planeringsfasen i medlemsstaterna och offentliggjorde riktlinjerna redan i juli 1999 , dvs. innan det nyvalda parlamentet hade inlett sitt arbete .
på det viset hindrade man parlamentet att påverka riktlinjernas utformning .
av den anledningen blir halvtidsbedömningen av artikel 42 i förordningen 1260 / 99 betydelsefull .
de nuvarande riktlinjerna utmärks generellt sett inte av klarhet och öppenhet .
trots att det är en viktig fråga berör de bara ytligt möjligheten att mäta de framsteg som gjorts utifrån verifierbara mål och i enlighet med gemenskapspolitikens strategier , och man uppehåller sig inte i tillräckligt hög grad vid utvidgningens effekter , och inte heller innehåller riktlinjerna specifika föreskrifter eller förtydliganden i frågan , vare sig för de regionala och nationella myndigheterna eller för kandidatländerna .
men oavsett detta är vi trots allt positiva till att man i riktlinjerna ställer de geografiska målen åt sidan och riktar in sig på sektoriell politik .
även om detta , teoretiskt sett , kan uppfylla kravet på koncentration och därmed kravet att åtgärderna skall vara effektiva , så uppkommer spontant frågan om den nuvarande situationen i mål 1-området är sådan att den faktiskt gör en integrerad politik möjlig . för att fullfölja en sådan skulle det krävas ett operativt samordnande instrument för avsättningarna .
vi kan därför , i princip , ge ett positivt svar på kommissionens begäran att få inrätta ett centrum för att främja strukturen i medlemsstaterna , men enbart genom att samordna förverkligandet och genomförandet av strukturella insatser på plats , så att ett sådant centrum inte blir till ett instrument för centralisering på övernationell nivå och att det garanterar att uppmärksamheten verkligen riktas mot de områden - jag säger det ännu en gång - som på grund av ett antal samverkande negativa faktorer ännu inte har nått upp till rätt nivå när det gäller att utnyttja strukturfonderna , för annars skulle det faktum att man ersätter det geografiska målet med sektorpolitik kunna sluta i en åtgärd som i själva verket blir negativ .
riktlinjerna innebär , i det skick de godkänts av kommissionen , en allvarlig begränsning eftersom de i stället för att uppfylla syftet att ange en inriktning räknar upp en katalog av tänkbara föreskrifter , en katalog som , eftersom den inte är prioriterad , i själva verket skulle kunna få medlemsstaterna att gå vilse genom att rikta deras uppmärksamhet mot ett brett urval av olika förslag , vilket skulle stå i strid mot den önskvärda koncentrationen .
vi skulle kunna säga att det verkar som om man ännu en gång har förlorat en chans att effektivt verka för en hållbar utveckling i städerna genom att bromsa den tilltagande urbaniseringen och den därmed följande förstöringen av landskapet .
man har inte i tillräckligt hög grad tagit hänsyn till betydelsen av generella subventioner , något som skulle kunna visa sig mycket användbart för att återskapa en balans mellan stad och land och dessutom vill man inte ge de lokala myndigheterna rätten att självständigt bestämma villkoren för en utveckling av sina territorier på kort sikt och genom egna åtgärder bidra till strukturfondernas reformansträngningar och till att målen effektivitet , koncentration och en snabbare byråkrati uppnås .
landsbygden måste äntligen betraktas som en tillgång som vi hela tiden måste investera mera i så att vi ger ungdomarna en anledning att stanna på landsbygden för att på så vis undvika att den faller sönder ekonomiskt och socialt .
det är ett numera välkänt faktum att för att uppnå det målet måste man i landsbygdsområdena skapa arbetstillfällen som inte bara är knutna till det traditionella jordbruket - även om det också är viktigt för att skydda miljön och den biologiska mångfalden - utan snarare inom sektorer som turism , idrott , kultur , miljö , små och medelstora företag , tjänster .
ett verkligt tomrum finns det i riktlinjerna på grund av bristen på konkreta förslag för att förverkliga samordningen mellan strukturfonderna och en strategi för ökad sysselsättning , en samordning som , just därför att den tillämpas för första gången under programperioden 2000-2006 , förutsätter att medlemsstaterna har behov av &quot; riktlinjer &quot; .
det bör även understrykas att kommissionen ännu en gång undviker problemet med konkreta åtgärder inom området lika möjligheter .
slutsatsen blir att detta är ett dokument som inte är särskilt tillfredsställande och i vissa avseenden en ren besvikelse .
betänkande ( a5-0107 / 1999 ) av berend
- ( pt ) vi stöder i det väsentliga den bedömning och de överväganden föredraganden gör angående den sjätte periodiska rapporten om den sociala och ekonomiska situationen och utvecklingen i europeiska unionens regioner .
vi begränsar oss därför till att betona några aspekter .
för det första , och som kommissionen själv säger , berodde de kraftiga framstegen i bni per capita i vissa fattiga regioner mellan 1991 och 1996 i hög grad på att de nya tyska delstaterna togs med i beräkningarna av gemenskapens genomsnitt , från första året , vilket var uppenbart avgörande för den påtagliga minskningen av unionens bni per capita .
därefter anser vi det vara av särskild betydelse att konstatera att återhämtningen som har skett i vissa regioner åtföljdes av en mycket liten ökning av sysselsättningen , något som därför kräver nya utvecklingsstrategier , med ett mycket större engagemang inom detta område .
denna situation talar emot en minskning av sysselsättningsskapande åtgärder till enbart medlemsstaterna , såsom föreslås i rapporten .
sist men inte minst , en hänvisning till föredragandens förslag om att denna typ av rapporter i framtiden , bland andra aspekter , också skall innehålla en analys av hur sammanhållningen mellan regioner i varje land utvecklas .
den mängd olika situationer och olika utvecklingsmönster som region för region uppvisas inom samma land , kräver i själva verket en fördjupad analys av denna fråga som gör det möjligt att förändra regionalpolitiken ( eller andra politikområden ) för att garantera sammanhållningen också inom varje medlemsstat .
berendbetänkandet erbjuder oss en intressant analys av den ekonomiska situationen och utvecklingen i europeiska unionens regioner .
men den franska delegationen i gruppen unionen för nationernas europa tar avstånd från vissa av de påståenden som finns i betänkandet .
punkt 26 &quot; påpekar att det särskilt behövs en konsolidering av budgeten såsom förutsättning för att den ekonomiska och monetära unionen och utvidgningen av unionen skall kunna genomföras med framgång &quot; .
när medlemsstaterna är förpliktade att genomgå en strikt finansiell bantningskur för att uppfylla konvergenskriterierna - det var för övrigt berättigat att de själva ansträngde sig för det - ger federalisterna prov på en mycket förvånande ekonomisk glupskhet .
för att visa att man erkänner emu : s och sammanhållningspolitikens misslyckande , säger man att bristen på uppnådda resultat beror på en brist på pengar . alla tävlar vältaligt om att kräva mer medel , men det finns ingen som funderar på om de utbetalade pengarna är effektiva .
vad skall man säga om ett budgetförfarande som går ut på att fastställa utgiftsmål i stället för utgiftstak , att - kosta vad det kosta vill - söka efter projekt för att med alla krafter spendera de anslagna medlen , i stället för att bevilja medel till befintliga projekt ?
utgiften blir ett mål i sig och ett bevis på att ett program har lyckats .
den statistik som europeiska kommissionen offentliggör i sin sjätte översikt visar trots allt , vilket berend underströk , den förda politikens begränsningar .
europeiska unionens rikaste regioner har ökat i betydelse mellan 1986 och 1996 , vilket vittnar om att rikedomar , arbetstillfällen och aktiviteter har koncentrerats till vissa områden : hamburg , bryssel , anvers , luxemburg , ile-de-france , darmstadt , oberbayern , bremen , wien , karlsruhe och emilia-romagna .
i motsats till vad föredraganden hävdar , kommer ekonomiska och monetära unionen att bidra till flykten från de mest avlägsna , mest lantliga och minst befolkade regionerna , till förmån för unionens centrala linje ( benelux , nordvästra tyskland , norditalien , île-de-france ... ) .
de fattigaste regionerna kommer steg för steg i kapp utvecklingsmässigt .
genomsnittet för de tio fattigaste regionerna uppnådde 41 procent av gemenskapens bnp år 1986 .
år 1996 låg det på 50 procent .
framstegen är särskilt tydliga i portugal och irland .
om de rikare blir allt rikare och de mycket fattiga blir mindre fattiga , verkar det som om genomsnittsregionerna , de som lyder under mål 2 , i realiteten har fått en lägre bnp , i vissa fall en icke försumbar minskning , samt försämrade sysselsättningsförhållanden .
det är särskilt tydligt i frankrike : i regionen champagne-ardennes , som jag har den äran att företräda , har bnp minskat från 105 till 94 procent av eu-genomsnittet , i pays-de-loire har den sjunkit från 95 till 91 procent , i auvergne från 89 till 83 procent .
detta är en generell tendens , som varken besparar rhône-alpes eller alsace .
den bekräftas i sverige och finland , länder där arbetslösheten under de senaste åren har ökat i oroande proportioner , liksom i flera av förenade kungarikets regioner .
därför kan det tyckas märkligt att mål 2 - vilket anslås till industri- och landsbygdsregioner som genomgår en ekonomisk omstrukturering - offrades i reformen av strukturfonderna till förmån för mål 1 och 3 : för perioden 1999-2006 ligger dess totalanslag på 22,5 miljarder ecu , en siffra som i princip är densamma som för perioden 1994-1999 .
de landsbygdsregioner som är berättigade till mål 5b kan räknas till de främsta offren för denna situation : i frankrike kommer 27 procent av den befolkning som är berättigade till strukturfonder att förlora sin rätt vid övergångsperiodens slut . denna siffra är mycket högre i vissa regioner , såsom pays de la loire , alsace och basse-normandie , högerns väljarbastioner som fallit offer för den pluralistiska vänsterregeringens politiskt förslagna klientilism .
med stöd av sådana beslut är det tveksamt om regionalpolitiken kan bidra till en harmonisk fysisk planering i europeiska unionens medlemsstater .
betänkande ( a5-0069 / 1999 ) av von wogau
med hänsyn till sysselsättningsläget i gemenskapen och europeiska unionens uttalade ambition att resolut bekämpa arbetslösheten , bör kommissionens analys av koncentrationer ta hänsyn till andra faktorer än konkurrensen .
som ett exempel skall jag ta upp företaget abb-alsthom power , som har en stor delegation anställda från hela europa närvarande i dag i strasbourg .
ledningen i abb-alsthom power , ett resultat av en fusion som genomfördes i juni 1999 , har tillkännagivit en omstrukturering som redan nu innebär att arbetstillfällen kommer att avvecklas i ett antal länder .
denna ödesdigra situation för sysselsättningen föranleder flera frågor , bl.a. om vilken information som har tillhandahållits det europeiska företagsrådet , som har funnits sedan 1996 .
och det förutsätter en förnyelse och förstärkning av gemenskapens direktiv om europeiska företagsråd .
det förutsätter också en kontroll av koncentrationer , vilken skall ta hänsyn till sysselsättningen , miljön och konsumenterna .
eftersom betänkandet från utskottet för ekonomi och valutafrågor är otillräckligt ur den synvinkeln , har jag avstått från att rösta .
- ( pt ) när kommissionen försöker tillämpa subsidiaritetsprincipen på gemenskapens konkurrenspolitik , decentraliserar man ansvaret för beslut och missbruk av dominerande ställning vad gäller företagsavtal som skapar snedvridning på marknaden , till nationella myndigheter och domstolar även om de fortfarande hör till anmälningssystemet för frågor om företagskoncentration och statligt stöd .
den ståndpunkt som nu har intagits är en strävan att skapa snabbare och billigare former för tillämpningen av konkurrenspolitiken , genom att eg-rätten tillämpas av de nationella domstolarna och inte av eg-domstolen , och även en inriktning mot specialdomstolar .
denna partiella åternationalisering av konkurrenspolitiken kan medföra ökade kostnader för medlemsstaterna .
å andra sidan , vilket föredraganden erinrar om , har ofta statliga monopol , i konkurrenspolitikens namn bytts ut mot privata monopol med privatisering av viktiga statliga sektorer och företag , så som är fallet i portugal , med negativa följder för landet och för dess arbetare .
kommissionens vitbok om en modernisering av reglerna om tillämpning av artiklarna 85 och 86 i eg-fördraget ( de nya 81 och 82 ) föreslår självklart inte en &quot; åternationalisering &quot; av konkurrenspolitiken , vilket vissa i europaparlamentet fruktar .
men den låter ana ganska intressanta utvecklingsmöjligheter för europeiska unionen .
kommissionen konstaterar att dess enheter översvämmas av förhandsanmälningar om avtal mellan företag som skulle kunna snedvrida konkurrensen , och fruktar att de kommer att bli fler när nya medlemmar tillkommer . den föreslår därför att man avskaffar det nuvarande systemet , dvs. att dessa avtal skall godkännas i förväg , och att tillämpningen av konkurrensreglerna skall decentraliseras till medlemsstatsnivå .
det mest anmärkningsvärda är enligt min mening den signal som detta förslag ger oss : kommissionen föregriper utvidgningens konsekvenser och anser att den med nödvändighet , ja nästan med automatik , förutsätter en reform av det centraliserade systemet .
denna reform består givetvis i en uppmjukning och inte en nedmontering .
på papperet skall kommissionen behålla kontrollen och den centrala ledningen i det nya systemet .
betänkandet av von wogau , som europaparlamentet just har röstat igenom , uppmuntrar för övrigt kommissionen på den punkten .
men samtidigt kan man lätt se att det sammanbrott som utvidgningen medför kan leda till en begränsning av gemenskapens behörigheter , och till en utvidgad subsidiaritet .
det är ett annat europa som på sikt kan komma att ta form .
är det förresten inte just det som skrämmer vissa socialister i europaparlamentet ?
de tyska socialdemokraterna röstade emot betänkandet av von wogau , eftersom de anser att det skulle sönderdela den europeiska konkurrenspolitiken , i klartext skada den likriktande överstaten .
märkligt nog har ett arbetsgivarparti anslutit sig till dem , eftersom det föredrar det europeiska systemet med &quot; en enda lucka &quot; , vilket för dem verkar vara mer ekonomiskt och mer stabilt juridiskt sett .
det är faktiskt en fördel med det nuvarande systemet .
men ur en annan synvinkel bör man också betänka att starten av den decentralisering som inleds i dag på sikt kan leda till en större frihet när det gäller hänsynstagandet till varje lands behov , något som kommer alla till del .
betänkande ( a5-0078 / 1999 ) av rapkay
de förtroendevalda i lutte ouvrière kommer inte att rösta för dessa betänkanden om den europeiska konkurrenspolitiken .
konkurrensen , dvs. det krig som de stora företagen för sinsemellan , tar sig ständigt uttryck i uppsägningar , nedläggningar av företag , för att inte tala om ett oändligt slöseri när det gäller utnyttjandet av den produktiva kapaciteten .
vi har fått ytterligare ett exempel på detta i och med att trusten abb alsthom power kommer att avveckla arbetstillfällen i europa .
18 miljoner arbetslösa , 50 miljoner fattiga i europeiska unionen , som trots allt är en av de rikaste regionerna i världen : däri ser vi resultatet av den konkurrens som eu-institutionerna har för avsikt att främja .
kommissionens vilja att reglera konkurrensvillkoren på den europeiska marknaden är löjeväckande , för den enda lag som konkurrensen lyder under är djungelns lag , dvs. att de mäktigaste krossar eller slukar de svagaste .
det är upprörande , framför allt ur en social synvinkel .
europeiska kommissionens rapport visar utan omsvep att unionens institutioner endast intresserar sig för de stora kapitalistiska företagsgrupperna , som hänger sig åt detta ekonomiska krig och inte på något sätt åt de offer som de själva skapar .
ingenting för att förhindra arbetslöshetens utbredning , ingenting för att skydda löntagarna , ingenting för att förhindra att de stora företagen driver en del av befolkningen till armod enbart för att skapa ännu större rikedomar för sina aktieägare !
skall vi medge att det finns en fördel med denna rapport , är det att den visar för samhällets arbetande majoritet att den inte kan hoppas på att eu-institutionerna kommer att upprätthålla , och än mindre förbättra deras levnadsvillkor .
genom att rösta emot detta betänkande gör vi oss till talesmän för alla dem som , i seattle och överallt i europa , har markerat sitt motstånd till en värld som reduceras till en strikt handelslogik .
vi röstar mot detta betänkande med omsorg om utvecklingen av de allmännyttiga tjänsterna , och i synnerhet till minne av offren för tågolyckan i paddington . deras död var inte ett olycksöde utan berodde på en absurd iver att konkurrensutsätta det som borde regleras .
detta betänkande är i grunden en lågt stående text , som endast inspireras av djungelns lag , för konkurrens kan inte lösa något av de problem som mänskligheten står inför vid detta sekelskifte .
vare sig det handlar om balansen i biosfären , att främja kulturen eller samarbeta med tredje världen , är en överdriven konkurrens en faktor som hänger samman med tillbakagång och osäkerhet .
och de 18 miljoner arbetslösa i europa , tror ni att de är offer för en alltför blygsam tillämpning av konkurrenspolitiken ?
vi är övertygade om motsatsen , och vi anser inte heller att de statliga stöden per definition är för stora .
enligt vilken dogm eller vilka effektivitetskriterier skulle de vara för stora ?
anser ni slutligen att det efter seattle är seriöst att förespråka en utvidgad roll för wto ?
endast de multinationella bolagens juridiska rådgivare kan ge prov på en sådan envishet .
betänkande ( a5-0087 / 1999 ) av jonckheer
jag gläder mig åt kvaliteten på den sjunde översikten över statliga stöd i eu och att den numera publiceras årligen , samt åt det faktum att generaldirektoratet för konkurrens använder sin webbplats för att ge både övergripande och mer detaljerad information till allmänheten .
jag tycker att föredraganden har en bra syn på statliga stöd , och jag vill gratulera honom till det .
man tenderar alltför ofta att sammanblanda statliga stöd med åtgärder som snedvrider konkurrensen .
visserligen är en effektiv konkurrenspolitik en förutsättning för att den inre marknaden och den ekonomiska och monetära unionen skall fungera väl .
samtidigt är den här typen av stöd ibland nödvändiga , vilket föredraganden betonar , och bidrar inte bara till att särskilda företag kan överleva , utan också till en hållbar utveckling ( artikel 6 i fördraget ) , tjänster av allmänt intresse ( artikel 16 ) samt ekonomisk och social sammanhållning ( artikel 158 ) .
det är likväl uppenbart att stöden måste kontrolleras , ett uppdrag som åligger europeiska kommissionen .
de stöd som unionens medlemsstater varje år anslår till de granskade sektorerna uppgick till totalt 95 miljarder euro under perioden 1995-1997 , varav 40 procent till tillverkningssektorn .
det är en avsevärd minskning i förhållande till den föregående perioden , 1993-1995 ( en minskning på 13 procent av det totala beloppet och en minskning från 3,8 till 2,6 procent av stöden till tillverkningssektorn ) .
de minskade stöden kan huvudsakligen förklaras med att stöden till tysklands nya &quot; länder &quot; har gått tillbaka .
i likhet med föredraganden beklagar jag att de siffror som presenteras i översikten inte täcker samtliga former av statliga stöd .
europeiska kommissionen bör snarast komma tillrätta med dessa brister .
den bör också samarbeta med medlemsstaterna för att i god tid förbättra kvaliteten på uppgifterna , dvs. inför den nionde översikten .
det vore bra om kommissionen offentliggjorde ett register som omfattar beloppen för statliga stöd per medlemsstat .
jag beklagar också att europaparlamentet är helt utestängt från den rådgivande kommittén om statliga stöd .
för att kompensera detta bör europeiska kommissionen lägga fram regelbundna rapporter för oss .
jag skall avsluta om en aspekt av utnyttjande av statliga stöd som jag tycker verkar särskilt farlig : det gäller de stöd som leder till omlokaliseringar av företag från en medlemsstat till en annan , vilket riskerar att skapa en jakt på subventioner som inte tillför eu : s gemensamma mål någonting .
därför skulle jag önska att nästa rapport om statliga stöd innehåller en utvärdering av statsstödens effekter på sysselsättningen och mottagarländernas industri och hantverk .
betänkande ( a5-0073 / 1999 ) av langen
i den viktiga konkurrensdebatten uttalade jag mig i förmiddags om langens text , som gäller tillämpningen av den sjätte regeln för stöd till stålsektorn under 1998 .
precis som eg-domstolen slog fast i beslut av den 3 maj 1996 är stålsektorn särskilt känslig för konkurrensrelaterade störningar .
därför var det berättigat att inrätta ett stödsystem för denna sektor , med ändamålet att garantera de livsdugliga företagens överlevnad , trots att artikel 4 c i eksg-fördraget förbjuder alla former av statliga stöd till stålsektorn .
detta är själva syftet med den sjätte regeln om stöd till stålindustrin .
samtidigt är det givetvis viktigt att förhindra att konkurrensvillkoren kränks och att marknaderna utsätts för allvarliga störningar , varför den här typen av stöd måste regleras .
det är således nödvändigt att även i fortsättningen begränsa de statliga stöden till att avse forskning , utveckling , miljöskydd samt stöd i händelse av företagsnedläggningar .
på samma sätt är det ytterst viktigt att medlemsstaterna uppfyller sin förpliktelse att till kommissionen anmäla vilka stöd som beviljats deras stålföretag , vilket artikel 7 i de aktuella reglerna föreskriver .
kommissionen föreslår att staterna skall sända in rapporterna inom två månader efter varje halvårsskifte , och under alla omständigheter en gång per år , utan att kommissionen skall behöva påminna dem om detta .
i likhet med föredraganden gladde jag mig åt kommissionens rapport , men jag beklagade att den inte täcker alla aspekter av statliga stöd .
även om reglerna för stöd till stålsektorn formuleras på ett mycket tydligt sätt , har kommissionen vid ett flertal tillfällen godkänt stöd till stålföretag som inte tillhör de kategorier som åsyftas i reglerna .
med omsorg om jämlikhet borde reglerna för statsstöd antingen tillämpas strikt eller ändras , om kommissionen vill godkänna andra stöd än dem som just nu är rättsligt tillåtna .
slutligen problemet med att eksg-fördraget löper ut .
stödsystemet bör finnas kvar efter år 2002 .
på denna punkt är det min uppfattning att endast en förordning från rådet kan ge erforderlig rättslig säkerhet och garantera ett formellt förbud mot alla de stöd som inte täcks av gemenskapens regler .
av alla dessa skäl har jag röstat för langenbetänkandet , och jag förväntar mig nu att kommissionen bemöter våra förfrågningar och krav .
oljebälte vid franska kusten
nästa punkt på föredragningslistan är kommissionens uttalande om oljebältet vid franska kusten .
härmed överlämnar jag ordet till kommissionens företrädare de palacio , som får inleda debatten .
herr talman ! jag uttalar mig å ppe-gruppens vägnar , men också i egenskap av förtroendevald från bretagne som är direkt berörd och chockad av dessa händelser .
tillsammans med franoise grosstête och ppe har vi ingivit ett resolutionsförslag .
i dag har vi ett kompromissförslag framför oss , vilket gläder mig .
erikas haveri är en europeisk angelägenhet , dels för att det förvanskar och smutsar ned några av europas vackraste stränder , med mycket allvarliga konsekvenser för turismen , dem som har havet som sin utkomst och de som försvarar miljön , och dels för att detta handlar om regler och kontroller som naturligt sett bör vara europeiska .
en katastrof som denna skulle i princip inte ha kunnat inträffa utanför de amerikanska kusterna . varför ?
därför att amerikanerna har tagit lärdom av exxon valdez-katastrofen och därför att de år 1990 utarbetade oil pollution act . denna akt utkräver ett större ansvar då den kan göra befraktaren ansvarig , den är dessutom mer tvingande och framför allt bättre kontrollerad genom en rad förordningar och i synnerhet den amerikanska kustbevakningen .
hade vi haft sådana bestämmelser , jag upprepar detta , hade katastrofen utan tvivel aldrig inträffat .
därför anser jag att vi måste se över de tillämpliga texterna , och särskilt det protokoll från 1992 som fråntog befraktarna allt ansvar , i det här fallet oljebefraktaren .
om befraktaren inte är ansvarig blandar han sig givetvis mindre i de kontroller som ligger på oljebolagens ansvar .
vi måste således se över bestämmelserna , och jag tackar er , fru kommissionär , för att ni pekade på alla de nuvarande bristerna i de europeiska bestämmelserna .
i övrigt krävs det , vilket ni nämnde , framför allt förstärkta kontroller - de kontroller som utförs av den stat under vars flagg fartyget seglar och de som utförs av klassificeringssällskapen .
ni sade att rina var ett italienskt klassificeringsregister som har godkänts av kommissionen .
på vilka grunder ges detta godkännande ?
vilka är garantierna om driftsäkerhet ?
ni kommer att sända en delegation .
vi väntar på resultaten med stort intresse .
man bör också stärka kustmyndigheternas kontroll och kontrollen i europeiska hamnar .
man skall komma ihåg att det finns en skrivelse från paris som förutsätter en minimikontroll : en fjärdedel av de båtar som lägger ut från en europeisk hamn måste kontrolleras av det berörda landets kustmyndigheter .
denna förpliktelse respekteras inte , varken i frankrike eller i många andra europeiska länder .
frågan är bara vilka konsekvenser kommissionen redan har tagit eller är beredd att ta ?
det förefaller också nödvändigt att förstärka den kontroll som befraktaren ansvarar för , i det här fallet oljebolaget .
om det har ett finansiellt ansvar , kommer denna kontroll utan tvivel att bli bättre .
till sist krävs det en samordning mellan olika kustmyndigheter för att nå fram till en europeisk gruppering , i likhet med de kustvakter som övervakar förenta staternas kuster .
herr talman ! varje gång en sådan här katastrof inträffar säger man att det aldrig får hända igen .
i verkligheten kan vi aldrig sätta stopp för olyckor till havs , men det åligger oss alla att dra lärdom när en sådan här olycka inträffar och använda denna lärdom för att minska riskerna i framtiden .
erika-olyckan var allvarlig , särskilt för de människor i bretagne som påverkas närmast , men den var förödande för stora delar av europas djurliv .
vissa säger att det var den värsta olycka som någonsin har drabbat fågellivet i denna del av europa .
det brittiska kungliga fågelskyddssällskapet tror att så många som 400 000 fåglar , kanske mestadels alkor , kan ha dött .
de bilder många av oss har sett på oljeindränkta fåglar som avlivas av veterinärpersonal var både sorgliga och tragiska .
vi vill alla ha högsta möjliga standard på fartyg oberoende av vilken flagg de för .
vi måste kräva efterlevnad av reglerna och se till att principen om att den som förorenar skall betala tillämpas så att ekonomiska straff och vissa incitament används för att sätta press på både rederier och oljebolag så att en bästa praxis införs .
jag instämmer i vartenda ord kommissionären sade i sina kommentarer , men frågan är hur lång tid det kommer att ta att tillse att åtgärder genomförs för att ta itu med problemet på det sätt hon föreslår ?
som politiker måste hon påminna sina tjänstemän om hur svårt det skulle bli om hon skulle behöva komma tillbaka till detta parlament om ett år om en liknande , precis lika förödande olycka skulle inträffa , och vissa av de åtgärder hon föreslår i dag fortfarande bara vore vackra ord som hon inte hade haft möjlighet att omsätta i verklighet .
tanken på att en olycka av detta slag kan inträffa inom en nära framtid bör bidra till att skärpa hennes och hennes tjänstemäns sinnen på ett fantastiskt sätt .
jag har tagit med en liten present till er : det är en oljekoka som en invånare på ön noirmoutier har skickat till mig , och hon skriver följande : &quot; varje gång det är flod täcks stranden av tung olja som läckt från erika .
varje gång det är flod tar frivilliga , militärer och brandmän fram enorma kokor av denna svarta klibbiga och tjocka tjära .
när blir det rent igen , när blir det ett slut på denna ödesdigra olycka ? &quot;
ja erikas haveri , liksom den ryska båtens haveri i turkiet för övrigt , kan inte accepteras eller tolereras med tanke på att den tekniska utvecklingen står på sin höjdpunkt .
det är dessutom oacceptabelt om man betänker att olyckan inträffade 20 år efter amoko cadiz-katastrofen , när man redan har sagt och flera gånger upprepat : &quot; aldrig mer ! &quot;
det är självklart politikernas , och därmed vårt ansvar att garantera säkerheten vid transporter till havs .
vi måste verkligen försäkra medborgarna att en liknande olycka aldrig mer kommer att inträffa .
men vi blir något frustrerade när vi lyssnar till er , fru kommissionär , för de som redan har ägnat sig åt den här typen av frågor vet att kommissionen och parlamentet förberedde , jag tror det var 1992 , en mycket intressant text , som redan då innehöll alla de förslag som finns i dagens resolution från utskottet för regionalpolitik , transport och turism .
det måste upprepas och upprepas igen : erika var en katastrof för mycket .
därför är det brådskande att europeiska unionen inleder en genomgripande revidering av direktiven om transporter till havs , för att göra dem mer tvingande samt upprättar en klar och detaljerad ansvarsordning för lastens ägare .
man bör t.ex. känna till att såväl shell som british petroleum vägrade att använda erika för sina oljetransporter .
varför medger man inte under dessa omständigheter att befraktaren , total , har ett ansvar ?
i era förslag bör ni även kräva dubbla fartygsskrov och att förbudet mot tankrengöring till havs verkligen respekteras .
man måste inrätta en europeisk inspektörskår , så att de verkligen och effektivt kan kontrollera båtarnas skick .
det är för övrigt lika brådskande att europeiska unionen åtar sig att reformera internationella sjöfartsorganisationen ( imo ) .
för vad tjänar det till att utarbeta bindande direktiv , om sedan flertalet båtar gör vad de vill när de väl är ute till havs ?
till sist , mina damer och herrar , vill jag skänka en öm tanke till alla frivilliga , natur- och fågelvänner , som spontant och generöst har anmält sig för att rädda oljeindränkta fåglar , genom att organisera en räddning med de medel som står till förfogande .
jag kan intyga att det är ett anmärkningsvärt arbete .
ni känner utan tvivel till att omkring 200 000 fåglar kommer att gå under i detta oljebälte , som är en oerhörd miljökatastrof och som praktiskt taget saknar tidigare motsvarighet .
ni vet också hur svårt det är i dag att bevara djurarter och hur svårt det är att bevara naturområden .
på den punkten , fru kommissionär , sade ni ingenting , dvs. hur kommissionen avser att bidra till återställandet av naturen och livsmiljöerna .
än en gång kommer ingen ansvarig att utpekas klart och tydligt .
i väntan på det är det alltid naturen som tar stryk .
herr talman ! min grupp begärde denna debatt för att ge parlamentet tillfälle att uttrycka sin solidaritet med de personer som är direkt berörda av miljökatastrofen , såväl i sin ekonomiska verksamhet som sina känslomässiga relationer med naturen .
tillåt mig att välkomna talesmannen för kollektivet &quot; oljebältet &quot; , bestående av medborgare från departementet morbihan ; javette-le besque , som har tagit plats på åhörarläktaren .
att uttrycka sin solidaritet , det har många frivilliga från frankrike och olika europeiska länder gjort genom att ge en viktig hjälpande hand till de drabbade .
att uttrycka vår , europaparlamentets solidaritet , det är i första hand att agera för att omedelbart få fram ett katastrofstöd till de familjer som drabbats av oljebältet . det innebär också att kräva en kvalitativ förstärkning av europeiska och internationella regler och säkerhetsnormer för transporter till havs , med tätare kontroller och mycket mer avskräckande sanktioner gentemot dem som bryter mot reglerna .
våra förslag avser bl.a. oljetankrarnas ålder .
bland dem som kontrollerades och bedömdes som bristfälliga förra året , var 15 av dem 20 år eller äldre , vissa mer än 30 och t.o.m. ännu äldre .
vidare bekvämlighetsflaggade fartyg .
enligt internationella transportfederationen seglade 40 procent av de fartyg som havererade 1998 under bekvämlighetsflagg , en symbol för vinst och utnyttjande av människor till förfång för säkerheten .
slutligen bristen på öppenhet .
man gör allt för att mörklägga kedjan av ansvariga , ägarnas identitet och de verkliga beslutsfattarna .
i alla dessa avseenden måste vi utverka verkliga och betydelsefulla förändringar , bl.a. en tidsfrist för inrättandet av nya normer som dubbla fartygsskrov . de som inte uppfyller kraven skall inte få lägga ut från hamnarna eller kryssa på medlemsstaternas vatten .
vi måste också uppnå ytterst strikta regler när det gäller utfärdande av sjövärdighetscertifikat och bedömningen av fartygens skick och underhåll .
vi måste slutligen se till att alla som bär ansvaret för en katastrof också bidrar till reparationerna .
i det här fallet tänker jag på gruppen total-fina .
herr talman ! denna strategi kan europeiska unionen utveckla visavi internationella sjöfartsorganisationen .
då kommer vi att ha visat allmänheten att vi gör någon nytta , för den här gången väntar man sig tydlig och konkret handling .
herr talman , fru kommissionär ! i egenskap av förtroendevald från den franska atlantkusten , från vendée , vill jag först och främst uttrycka den upprördhet som offren för erikas oljebälte känner inför katastrofen , en katastrof som har förorsakats av - inte en naturkatastrof som de orkaner vi nyligen drabbades av - utan av en brottslig handling .
i det akuta läget och inför en stor prövning , uttrycktes en fantastisk solidaritet : en lokal solidaritet , en nationell solidaritet , en mellanstatlig solidaritet .
förväntningarna hos de drabbade befolkningarna , de som har förlorat allt - särskilt de som är yrkesmässigt beroende av havet och turismen - de vilkas verksamhet är ruinerad för flera år framöver , är inte bara att förorenarna skall betala för de skador de har åsamkat , utan också att man gör allt för att deras olycka skall hjälpa andra i framtiden och förhindra att liknande brott begås igen .
vi betalar givetvis priset för våra försummelser .
staterna gjorde nämligen bedömningen - med gemenskapens välsignelse - att det inte längre var lönsamt att ha en egen handelsflotta och lät därmed ett stort kunnande i skeppsbyggnad försvinna . därför kan vi inte längre spåra fartygens ursprung och därför får vi se riktiga vrak segla på våra farvatten under bekvämlighetsflagg , till förmån för de multinationella bolagens kortsiktiga intressen .
vi måste verkligen sätta stopp för denna ström av oansvarighet , oansvariga befraktare , skeppsredare som är omöjliga att hitta och eftergivna certifieringssällskap .
dagens läge är mycket förvirrat .
dessa frågor bör självklart hanteras på internationell nivå , men imo : s nuvarande internationella regler är otillräckliga och alltför släpphänta . varken medlemsländerna eller gemenskapen har varit påstridiga och försökt få till stånd striktare regler , trots tidigare inträffade katastrofer .
visserligen existerar internationella fonden mot oljeföroreningar ( fipol ) , men den sprider ut ansvaret och har alltför begränsade ramar , som därför måste ses över .
man bör absolut se över frågan om bekvämlighetsflagg inom ramen för imo .
det är medlemsstaternas och gemenskapens sak att vidta erforderliga åtgärder för det ändamålet .
jag vill erinra om att erika bekvämlighetsflaggades av en stat som har ansökt om medlemskap i unionen .
vi har också gemenskapens direktiv , men de tillämpas i ringa utsträckning eller inte alls , på grund av att de nationella kontrollanterna är alltför få .
vi måste snarast åtgärda den bristen .
ett direktiv om säkerhet till havs har förberetts under många år , men arbetet framskrider mycket långsamt .
på den punkten visar kommissionen en tröghet som inte kan tillåtas och en oförmåga som inte kan accepteras .
presentationen av kommissionens meddelande om denna centrala fråga skjuts ständigt upp och är nu planerad till juli , men den bör absolut tidigareläggas .
vad gäller de konkreta bestämmelserna måste de vara särskilt tydliga och strikta .
jag vill nämna tre som vår grupp prioriterar .
för det första måste tankerägarnas ansvar klart och tydligt fastställas , och de som faller offer för en förorening måste utan tvekan kunna ställa dem till svars .
det bästa sättet att förebygga olyckor inför framtiden , är att befraktarna kan vara förvissade om att de kommer att straffas hårt , civilrättsligt , straffrättsligt och finansiellt , om de inte är ytterst vaksamma beträffande säkerheten på de fartyg de väljer ut .
för det andra måste kravet på dubbla fartygsskrov för oljetankrar som får segla på gemenskapens farvatten införas så snart som möjligt , och inte uppskjutas på obestämd tid .
för det tredje måste man snarast fastställa en strikt begränsning av åldern på de fartyg som tillåts frekventera gemenskapens farvatten .
maximiåldern skulle kunna vara 15 år .
lyckas man inte uppnå en tillräckligt tydlig , strikt och rigorös ram på gemenskapsnivå , bör de medlemsstater som för egen del vill införa striktare bestämmelser tillåtas att göra det för att skydda sin befolkning och sitt territorium , på samma sätt som förenta staterna tog lärdom av exxon valdez-katastrofen genom att kräva dubbla fartygsskrov och förbjuda alla fartyg som är äldre än 20 år att segla på deras farvatten .
förenta staterna skulle således ha vägrat erika tillträde till sina farvatten .
om gemenskapen hade gjort detsamma hade en oerhörd katastrof kunnat undvikas .
herr talman , fru kommissionär ! låt oss denna gång verkligen ta lärdom , även när massmedias och parlamentsledamöternas känslor har lagt sig .
herr talman ! torrey canyon , olympic bravery , haven , amoko cadiz , gino , tanio ; detta är en rad namn som är förknippade med dystra minnen .
och nu erika .
vems tur är det sedan ? 21 år efter amoko cadiz får vi för femtielfte gången se ett oljebälte , det sjunde sedan 1967 och beviset för alla efterföljande regeringars oansvarighet .
västra atlanten får än en gång betala ett högt pris för deras oförmåga att reagera , för att de kapitulerar inför de multinationella bolagen .
det är svårt att förstå varför fransmännen och européerna tillåter det som amerikanerna förbjuder , och varför europa , som normalt sett är så snabbt på att lagstifta i miljöfrågor , inte har gjort något för säkerheten till havs .
resultatet ser vi i dag .
erika , ett fartyg som seglade under maltesisk flagg , ett flytande vrak som klassas som en av de farligaste oljetankrarna , har smutsat ned våra kuster längs en drygt 400 km lång sträcka , vilket är en långt mer allvarlig förorening än den som amoko cadiz förorsakade .
som förtroendevald från loire-atlantique kan jag tyvärr intyga det .
dessa upprepade katastrofer hänger på inte på något sätt samman med naturens krafter , det finns inget ödesbestämt över dem .
de är en konsekvens av människors inkonsekvens .
detta är en riktig miljökatastrof .
endast de som inte har varit där och sett den hårda verkligheten kan betvivla det .
det är också en ekonomisk katastrof för alla dem som lever av havet och turismen ; fiskare , ostronodlare , musselodlare , salinarbetare , handlare , osv.
svepeskålen erika måste bli den sista i raden .
vi måste först och främst göra allt för att bringa klarhet i haveriet .
varför inte utse en parlamentarisk undersökningskommitté eller låta parlamentsledamöter delta i den delegation som kommissionen aviserade för en stund sedan ?
sedan måste vi snarast anta lagar som fordrar grundligare kunskaper om det transporterade godsets egenskaper .
enligt experterna skulle oljan från erika ha sjunkit till bottnen och aldrig ha nått kusterna .
men vi vet vad som hände .
det krävs vidare att man inför en tillförlitlig teknisk kontroll , i likhet med frankrikes obligatoriska tekniska kontroll av fartyg som är äldre än fem år .
det krävs bestämmelser för användningen av bekvämlighetsflagg , krav på dubbla fartygsskrov för transporter av förorenande och farliga ämnen och en utveckling av tekniken för att hantera och samla upp oljeutsläpp .
det är enligt min mening ett minimum på tröskeln till det tredje årtusendet .
de fartyg som inte uppfyller kraven måste nekas tillträde till europeiska farvatten ; förorenarnas , skeppsredarnas och befraktarnas ansvar måste fastställas enligt principen &quot; den som förorenar skall betala &quot; ; övervakningen på haven måste förstärkas för att förhindra tankrengöring ; en seriös och tillförlitlig kontroll av fartygstankrarna måste införas ; en konsekvent budgetpost för &quot; naturkatastrofer &quot; måste återupprättas för medlemsländerna , och i väntan på det bör man uppbåda ett exceptionellt gemenskapsstöd och se till att medel ur strukturfonderna kan anslås till de katastrofdrabbade departementen .
å edd-gruppens vägnar har jag också ingivit en resolution i den frågan .
herr talman ! under de senaste åren har det över hela världen förekommit upprepade svåra katastrofer med tankfartyg , utan att några nämnvärda eller effektiva motåtgärder har vidtagits .
denna gång är det särskilt illa , inte minst därför att det har drabbat en stor europeisk stat , en händelse som kan upprepas när som helst .
för att minska dessa risker behöver vi snarast ett direktiv .
de 15 räcker uppenbarligen inte .
dessa garanterar - utan anspråk på att vara fullständiga - minst 3 punkter : inget skrotfärdigt tank- eller fraktfartyg får någonsin mer anlöpa en hamn i europeiska unionen .
alla inblandade , inklusive den som beordrat transporten , är ansvariga för följdskadorna , och tillräckliga försäkringar måste tecknas av dessa inblandade .
endast på så sätt kan de drabbade ha en chans att få sina skadeersättningsanspråk tillgodosedda .
men vi måste vara klara över att det långsiktiga målet måste sättas mycket högre .
det betyder att vi behöver en verklig kostnadsuppskattning för vårt hela energiförsörjningssystem .
herr talman ! skulle jag kunna få börja med att rikta ett stort tack till kommissionär palacio för det klara , adekvata och även mycket rakryggade svaret .
tusen tack för detta .
det innebär också att jag i varje fall har stor respekt för det briefing-pm som hon skickade den 10 januari , men också för de åtgärdspunkter som hon tillkännagav i dag .
katastrofen med erika visar att när övergripande trafik- och transportbestämmelser saknas på internationell och europeisk nivå så är det naturen och miljön som drar det kortaste strået .
den skada som har uppstått , även på det ekologiska området , går inte att uttrycka i pengar .
det är anledningen till denna gemensamma debatt med kollegerna från transport och miljö .
under julferien när de nederländska medierna uppmärksammade katastrofen med erika gick jag ut på internet för att se vilka åtgärder det nu egentligen var som skulle vidtas , i synnerhet efter det att premiärminister jospin hade sagt att europa måste göra mer .
vad jag förstod av detta var att det egentligen finns tillräcklig lagstiftning , men att problemet är att det inte sker några kontroller .
jag skulle här vilja uppmärksamma ett par punkter , som även kommissionären nämnt i förbigående .
först och främst port-state control , de 25 procent av alla fartyg som måste kontrolleras .
jag tror att dessa 25 procent inte bara måste upprätthållas , utan att man därefter också måste sörja för att det görs fler kontroller ; dessa 25 procent måste således höjas .
när ett skepp inte längre får segla måste inte bara sakförhållandena kontrolleras , utan det måste också inrättas ett rättsligt system där man säger : det är klokast att ni inte går ut till havs mer eller det får ni inte göra längre .
men något sådant finns inte .
herr talman ! på den punkten skulle jag gärna se att det hände något .
slutligen något om de tekniska krav som ställs på fartyg ; mina kolleger talade nyss om att det i förenta staterna sedan 1999 i varje fall måste finnas dubbla kölar .
jag anser att vi måste gå längre på den punkten , och jag anser också att marpol-fördraget , som träder i kraft 2001 , måste ses över ordentligt .
herr talman ! sedan måste man också kritiskt se över anslutningsförhandlingarna med malta , och jag vill framföra mitt tack och min beundran till de många icke-statliga organisationer som i varje fall har tagit upp händerna ur byxfickorna för att rädda djur .
herr talman ! vi har redan ofta fört denna diskussion .
vi har hittills inte uppnått någonting , och vi har inte kunnat enas här i europeiska unionen .
därför tror jag att det bara är meningsfullt med dagens debatt om det som vi alla säger i dag , och det som ni , fru kommissionär , här har tillkännagett , faktiskt utmynnar i en lagstiftning , dvs. om ni säger till alla era regeringschefer och era ministrar : detta måste ni genomdriva i ministerrådet .
låt mig på förhand säga att vi talar om en miljökatastrof , som också har ekonomiska effekter och hotar existenser .
vad måste vi nu göra ?
jag vill ju alls inte gå tillbaka till det förflutna . jag vill se framåt .
jag vill säga något om vad vi måste göra .
naturligtvis behöver vi fartyg med dubbelt skrov .
det är klart , men detta är något som bara kommer att få effekt på medellång och lång sikt .
vad behöver vi då genast ?
vi behöver en teknisk kontroll av fartygen , nämligen en bindande teknisk kontroll av fartygen vartannat år , och utan detta certifikat får inget fartyg framföras .
det behöver vi på europeisk nivå , och det behöver vi internationellt , som en teknisk övervakningsinstans , som en teknisk besiktning av fordon , vilken i tyskland måste göras vartannat år .
om man inte har något besiktningsinstrument , får man inte köra fordonet .
det behöver vi för fartyg .
för det tredje behöver vi en kontroll av dessa certifikat och ett försäkringsbevis i hamnarna , och detta i alla europeiska unionens hamnar .
om detta certifikat och försäkringsbevis saknas , beläggs fartyget med kvarstad och får trots alla hamnavgifter inte lämna hamnen .
där måste vi vara ense , i alla hamnar i europeiska unionen , från marseille via rotterdam till wilhelmshaven , cuxhaven och var än fartygen anlöper .
för det fjärde måste det finnas ett ansvar hos fartygsägaren , och inte bara skrattretande 12 miljoner dollar , utan minst 400 miljoner dollar , vilket han måste styrka med hjälp av försäkringsbevis .
då måste det finnas ett ansvar hos det land , under vars flagga fartyget seglar .
vi behöver den säkerheten att det land , under vars flagga fartyget seglar , i tveksamma fall övertar ansvaret .
det blir en underbar kontroll !
jag kan garantera att de länder som utdelar flaggorna då också kommer att se till att de inte måste bära ansvaret .
vi behöver för det femte den garantin att detta krävs för alla fartyg i europeiska unionens hamnar och farvatten , för övrigt också i kandidatländernas . det betyder att de krav som jag har nämnt gäller för alla farvatten .
slutligen behöver vi det allra viktigaste : vi behöver ha ett bra minne , ty vi kommer här under den närmaste tiden att oftare tala om lagstiftning .
vi kommer oftare att tala om miljönormer .
då vill jag inte att någon kommer och säger : dessa krav leder till att vi förlorar arbetstillfällen i hamnarna .
fackföreningarna kommer , industrin kommer .
vi behöver ett bra minne , kära kolleger .
här tittar jag på många av er , som hittills inte har gått i bräschen för miljörörelsen .
gå hem och säg : de normerna har vi hittills inte bekymrat oss om .
vi behöver ett bra minne när det gäller vad som krävs i hamnarna .
vi behöver ett bra minne , när vi säger : vi är ense vad beträffar hamnavgifter och hamnbestämmelser , och vi spelar inte ut den ena mot den andra i europeiska unionen .
om vi klarar av det , så kommer vi kanske om ett par år att ligga bättre till !
herr talman ! roth-behrendt uttryckte väldigt mycket av mina tankar .
vi har nu fått en perfekt uppräkning av olika åtgärder .
men hur använder vi det krismedvetande som denna ekologiska katastrof har lett till ?
jag jämför med när en tidigare generation införde plimsollmärket , en märkning som infördes för att undvika försäkringsbedrägerier med undermåliga fartyg .
var har vi samma krismedvetande som generationerna före oss hade ?
jag anser att det vi skall gå in för är den certifiering som roth-behrendt talar om , den märkning med gröna märken på tankfartyg som vissa hamnar i europa har fört på tal .
vi måste dessutom kritiskt granska klassificeringssällskapen .
jag tycker inte att vi kan acceptera deras förfarande .
vi behöver oberoende förfaranden och förfaranden med insyn .
slutligen vill jag säga att när mitt land ger miljöstöd till redare som vill förbättra miljökvaliteten , så finns det enheter inom kommissionen som betraktar detta som förbjudet varvsstöd .
den ena handen inom kommissionen vet inte vad den andra gör .
det är inget acceptabelt förfarande att man inte får göra miljöförbättrande åtgärder , som är i enlighet med kommissionens riktlinjer , eftersom dessa anses utgöra förbjudet varvsstöd .
herr talman ! vi kommer att rösta för resolutionen från gue / ngl-gruppen , eftersom den pekar ut total-fina som ansvarig för denna miljökatastrof , och eftersom jag skriver under på förslaget att förbjuda bekvämlighetsflagg och bruket av föråldrade båtar , och att införa ett krav på dubbla fartygsskrov för oljetankrar .
jag vill bara tillägga att det minsta man kan begära är att total betalar alla kostnader för de skador som oljebältet direkt och indirekt har förorsakat .
hur skall man kunna förhindra att liknande katastrofer inträffar igen om man inte vidtar ytterst stränga åtgärder gentemot de stora oljetrusterna , och även andra , som för att kamma in ytterligare vinster tar risken att göra vår planet obeboelig ?
hur är det möjligt att inte uppröras över att en bank vägrar lämna ut namnet på erikas ägare genom att hänvisa till banksekretessen , och att ingen regering reagerar på det ?
det egentliga problemet är att alla regeringar , liksom alla eu-institutioner , ger stora truster som total-fina och dess likar rätten att maximera vinsterna till nackdel för såväl sina anställda som miljön .
man tillerkänner företag och banker rätten att hemlighålla sina affärer , även om denna sekretess skyddar rent kriminella handlingar .
under dessa omständigheter kommer även de allra bästa resolutioner att förbli bevisningsfel , som inte kan förhindra att de stora trusterna åsamkar skador .
erika sjönk rakt framför mitt hem . hon ligger fortfarande där med 20 000 ton i sidorna , och man vet ännu inte vart dessa ton kommer att ta vägen .
hon hade kunnat sjunka någon annanstans .
men av en slump sjönk hon just där , och det bretagne som jag kommer ifrån skall inte behöva ursäkta sig för att det är en halvö , för bretagne får ofta uthärda skeppsbrott .
jag tänker framför allt på de 26 indiska sjömän som man inte talar om och som inte räddades .
människor hade kunnat dödats i den här katastrofen , och säkerhet till havs handlar främst om människoliv .
i dag är dessa sjömän ett avlägset minne .
det är ett mirakel om de har räddats .
så kommer man att börja om på nytt precis som för 20 år sedan med amoco , ett hugg på nordkusten , ett hugg på sydkusten , ett hugg på västkusten .
och det skulle kunna fortsätta på det viset .
fru kommissionär ! eftersom det är mycket ont om tid skulle jag bara vilja räkna upp de sju punkter som vi anser att det är ytterst viktigt att arbeta på , och ni har säkerligen nämnt några av dem : dubbla fartygsskrov så snart som möjligt på våra farvatten och en så strikt statlig kontroll som möjligt i hamnarna .
det krävs framför allt att klassificeringssällskapen är förpliktade att offentliggöra sina rapporter , eftersom de inte är kända .
vidare att de femton medlemsstaterna harmoniserar påföljderna - de får inte skilja sig åt , utan måste vara desamma överallt .
man måste skärpa bestämmelserna om bekvämlighetsflagg , inte för att de nödvändigtvis är sämre båtar , utan för att det finns många dåliga båtar som seglar under bekvämlighetsflagg ; förbättra informationen om samtliga fartyg i världen , vilket visserligen redan är planerat , och att ringa in och skärpa ansvaret .
i det avseendet skulle jag vilja veta vem som äger erika , för begreppet juridisk person i vår rätt är en sak , men det finns alltid fysiska personer bakom - var är de , erikas ägare ?
kanske i vackra villor vid vackra stränder för att sola sig .
vi skulle gärna se deras namn och deras ansikten .
och slutligen en förbättring av utbildningen för fartygsbesättningar .
i vårt samhälle finns det ingenting som en nollrisk , men vi kan åtminstone vara så försiktiga som möjligt .
herr talman ! jag välkomnar kommissionärens uttalande .
eftersom jag själv har tillbringat lång tid till sjöss är jag väl medveten om havets makt och destruktiva kraft som gör ändamålsenlig utformning och underhåll av skepp och båtar avgörande .
jag skulle vilja uttrycka mitt deltagande med alla dem som handskas med konsekvenserna av att oljetankern erika förliste och sjönk .
detta har varit en miljökatastrof liksom ett djupt beklagligt resursslöseri .
man bör notera att oljeindustrin , genom de internationella oljeskadefonderna , betraktar sig som ansvarig för över 90 procent av den beräknade kostnaden för denna olycka , eller cirka 170 miljoner dollar , enligt konventionen från 1969 och 1992 års protokoll .
detta tycker jag tyder på att vi också bör uppmana fartygens ägare , den stat vars flagg man för och kontrollmyndigheterna att ta sin del av ansvaret .
låt oss emellertid , innan vi rusar åstad med en hel räcka nya åtgärder och regler , noggrant titta på gällande bestämmelser så att vi är säkra på att de tillämpas på rätt sätt .
det är bättre att följa uppmaningar att modifiera och förbättra gällande lagstiftning än att inlåta sig på nya förslag .
i detta sammanhang stöder jag kraven på att utöka hamnkontrollen för att tillse att en total och effektiv kontroll görs .
jag stöder krav på att tillse att klassificeringssällskapen på ett effektivt sätt övervakar fartygens strukturella skick och hålls ansvariga för sina handlingar .
krav på förbättringar av skrovkonstruktionens utformning , speciellt fartyg med dubbla skrov , är förnuftiga men tar tid att genomföra i hela flottan .
det finns inget som kan ersätta rigorösa regelbundna kontroller .
herr talman ! jag vill framföra ett tack till mina socialistiska kolleger , i synnerhet till dem från utskottet för regionalpolitik , transport och turism samt utskottet för miljö , folkhälsa och konsumentfrågor , för att de inte har glömt att denna olycka även påverkar fiskerisektorn .
förutom skadorna på miljön , skadorna på ekosystemet som inte går att reparera och förlusterna för turistsektorn , innebär oljebältena ett dråpslag för fisket , för bevarandet av resurserna i havsmiljön , och det kommer att ta många år att återställa den förstörda kusten .
det är ingen tillfällighet , fru kommissionär , att de drabbade områdena alltid är europeiska regioner med en försenad utveckling , de regioner som hankar sig fram med hjälp av en kombination av turism och fiske , och där det i de flesta fall saknas andra resurser .
det är även dessa regioner , fru kommissionär , som under hela året får stå ut med vissa redares oförskämda agerande då de rengör botten på sina fartyg utanför kusten , utom all kontroll .
jag kommer själv från galicien , en region som tidigare har drabbats av liknande olyckor .
bretagne och galicien , två europeiska ändpunkter , blir ständigt offer för det bristande ansvarstagandet hos dem som väljer att bryta mot säkerhetsbestämmelserna och transportera råolja i fartyg som i sig utgör potentiella oljebälten .
därför anser jag att det är nödvändigt att agera i två olika avseenden .
för det första genom att vi ber att kommissionen , inom ramen för det planerade stödet till fiskerisektorn , vidtar särskilda åtgärder för att mildra effekterna av denna katastrof för den produktiva sektorn i de drabbade regionerna , och att vi dessutom ber kommissionen av sig själv och de internationella organen kräva en striktare kontroll av fartyg med bekvämlighetsflagg .
därför bör man under den pågående förhandlingsprocessen om maltas anslutning till europeiska unionen passa på att kräva att malta utövar en sträng kontroll av oljetankfartyg under deras flagg .
för det andra måste vi agera förebyggande .
portugal är ett land där man tydligt visat hur känslig man är för frågor med anknytning till havet .
jag skulle vilja uppmana det portugisiska ordförandeskapet att undersöka möjligheten att införa en övergripande strategi för att förebygga olyckor till sjöss på europeisk nivå , genom att man sammanför all de medel som står till vårt förfogande - tekniska , strukturella och socioekonomiska sådana - för att undvika en upprepning av en katastrof som denna i framtiden .
slutligen , herr talman , vill jag lyfta fram det arbete som har utförts av frivilliga och av de lokala myndigheterna , som påminner mig om gamla tider då jag - som borgmästarinna - fick uppleva liknande situationer .
vi måste tacka alla dem som i ett sådant utsatt läge med knappa resurser har visat mod i kampen mot de allvarliga konsekvenserna av denna katastrof för kustregionerna , ekosystemet till sjöss och europas fiskeresurser .
herr talman ! i egenskap av ordförande för utskottet för regionalpolitik och transport skulle jag vilja gratulera kommissionen , och speciellt kommissionsledamoten loyola de palacio , till deras sätt att hantera denna fråga , som har väckt så starka reaktioner i hela europa .
vi i transportutskottet är beredda att diskutera kommissionens meddelande om säkerhet till havs , och vi är naturligtvis också beredda att senare diskutera vilka konsekvenser detta meddelande får i rättsligt avseende .
sedan skulle jag vilja göra några påpekanden :
för det första ; det är med all rätt som kommissionen i sin undersökning framför allt söker utkräva ansvar av det italienska fartygsinspektionsbolaget rina , eftersom vi måste ta reda på om gemenskapsrätten har tillämpats .
detta bör vara utgångspunkten för våra ansträngningar .
för det andra ; förutom redarnas ansvar är det lämpligt att vi i sådana fall även beaktar befraktarnas ansvar , det gäller t.ex. oljebolagen som också bär ansvar för ekologiska katastrofer som i det här fallet , men som också måste ta sitt ansvar för att återställa det som skadats .
reaktionen på den ekologiska katastrofen är verkligen befogad .
men detta får inte leda till att vi skuldbelägger all handelssjöfart , som ju är en mycket viktig bransch för ekonomin , eftersom den svarar för ungefär 1 / 3 av transporterna , och därför bör våra reaktioner vara måttfulla , stränga men också korrekta .
jag motsätter mig inte alls att man överväger en skärpning av gemenskapsrätten men , såsom även andra kolleger har framhållit , vi bör utgå från tillämpningen , för det finns redan ett regelverk - och det får vi inte glömma - på europeiska unionens nivå .
detta regelverk är ganska avancerat - åtminstone om man jämför det med situationen på global nivå - och följaktligen är medlemsstaterna , under kommissionens överinseende , skyldiga att verkligen börja tillämpa gemenskapsrätten .
herr talman , fru kommissionär ! jag anser att den beklagansvärda händelsen med erika i själva verket , så som man har påpekat här i eftermiddag , bör bli en definitiv vändpunkt som markerar före och efter den här typen av olyckor i europeiska unionen , där det sedan 1967 har inträffat sjutton olyckor med stora oljetankfartyg , det vill säga mer än en olycka vartannat år .
de sociala och ekonomiska skadorna , som vi redan har talat om här i dag , både vad gäller en försämrad sysselsättning och försämrade resurser inom fiske och turism , är av den omfattningen att de mer än väl motiverar ett beslutsamt och övertygande agerande från gemenskapsinstitutionernas sida .
även jag , fru kommissionär , vill tacka för kommissionens snabba reaktion på denna händelse och de åtgärder man nu vidtar och de som är på gång .
och jag litar på att dessa åtgärder inom de närmaste månaderna leder fram till ett tydligt och övertygande rättsligt instrument - eventuellt ett direktiv - som en gång för alla sätter stopp för dessa pirater på 2000-talet , som berövar oss alla på havets rikedom och skönhet .
jag skulle vilja göra ett påpekande beträffande en av de åtgärder som kommer att vidtas och som har påtalats av kommissionären och av flera av mina kolleger .
det gäller dubbelskrovet , som innebär att lasten inte har kontakt med ytterskrovet , det vill säga skrovsidan mot sjön .
fru kommissionär , det finns många experter som anser att dubbelskrovet inte är tillräckligt säkert och i stället rekommenderar ett så kallat &quot; ekologiskt skrov &quot; , där havsvattnet vid en eventuell olycka tränger in i tankarna och gör att oljan , på grund av trycket , förs över till andra tankar .
jag anser , fru kommissionär , att det är dags att vi röstar på de säkraste tekniska åtgärder som finns .
därför anser jag att vi inte får nöja oss med att kopiera en lagstiftning som gäller i andra länder .
jag anser att vi kan och bör förbättra den lagstiftning som finns på området .
varje analys av kostnader och vinst där man beaktar de totala skadorna på människorna och miljön till följd av dessa olyckor , kommer att ge oss rätt .
jag skulle först och främst önska att vi gläder oss över vårt förfarande . det gör det möjligt för oss att slutligen lägga fram en gemensam resolution - efter det att alla politiska grupper har samlat sig för att uttrycka vad alla känner .
under dessa tragiska omständigheter tror jag att det vore en missuppfattning och en skam om vi talade med flera olika röster , principiellt sett .
det faktum att parlamentet i dag lägger fram en resolution med en enda röst - vi kunde konstatera de föregående talarnas samsyn - tror jag utgör ett tillfälle för oss parlamentariker att sätta press på ett antal regeringar , som tvekar och ägnar sig åt undanmanövrar , och jag tror att det är en mycket stark politisk handling som vi lägger i kommissionens händer för att förbereda ett europeiskt maritimt område .
jag tror att det står helt klart - och det är den första slutsatsen man kan dra av erikas katastrof - att allmänheten inte skulle förstå varför man antar bestämmelser för choklad men inte för transporter till havs .
allmänheten skulle inte förstå varför man talar om ett gemensamt rättsområde , att man talar om ett gemensamt luftområde , att man talar om ett gemensamt järnvägsområde och en gemensam marknad , men inte om ett maritimt område .
i dag tror jag att det är ett arbete som måste inledas med en bestämd vilja till resultat , konkreta resultat .
kommissionären pekade på tre stora avsnitt som bör utvecklas : en modernisering av vår lagstiftning , så att vi kan ta fram normer .
till min stora tillfredsställelse noterade jag för övrigt att t.o.m. de euroskeptiska grupperna , som förespråkar staternas suveränitet , vädjar till europa att fastställa bestämmelser , och jag tror att eu är rätt nivå för det .
ibland reglerar vi saker som i stor utsträckning skulle kunna regleras på en lägre nivå .
på det här området bör vi ge ett svar till allmänheten .
det är mycket viktigt och alla måste känna sig berörda , för när allt kommer omkring är vi internationellt sett inte mer än en halvö .
det krävs således uppföljningsregler .
efter en modernisering av vår lagstiftning måste vi också inrätta systematiska kontroller och slutligen tillämpa principen om förorenarens / den betalningsskyldiges ansvar , vilket självklart är en förebyggande princip .
jag skall strax avsluta , men jag vill också säga att jag har lämnat en förfrågan till utskottet för transport och turism om en offentlig utfrågning , för att vi direkt skall kunna följa upp ärendet erika och förse framtida reflektionsarbeten med nytt underlag .
jag hoppas att alla politiska grupper kommer att stödja vår förfrågan om en offentlig utfrågning .
herr talman ! oljetankern erika , vars ägandeförhållanden döljs av brevlådeföretag på malta och kanske italien och grekland , hyrd av totalfina för transport av olja , förliste utanför den bretagniska kusten med alla katastrofala följder det medfört .
konsekvenserna för miljön , den europeiska havsmiljöns flora och fauna är enorma .
orsaken till katastrofen måste sökas i oljetankerns försvagade struktur .
folk tvivlar således på säkerheten för fartyg som transporterar farlig eller förorenande last .
den internationella maritima organisationen har utgivit en internationell reglering för detta .
stater kan utföra hamninspektioner .
i europa är lagstiftningen strängare och man måste , är förpliktigad , att kontrollera 25 procent av de inlöpande fartygen enligt direktivet port-state control .
men det verkar som om inte en enda medlemsstat uppnår denna procentandel på grund av brist på inspektörer .
det står helt klart att det inte råder brist på lagstiftning .
jag tror att kommissionären har alldeles rätt i det .
det som fattas är tillämpning av den redan befintliga lagstiftningen .
men hur skall det nu gå till när vi faktiskt har brist på inspektörer , ärade europeiska kommission ?
kan kommissionen försäkra att direktiv 93 / 75 om minimikrav för fartyg som anlöper eller avgår från gemenskapens hamnar med farligt eller förorenande gods verkställs på ett korrekt sätt i alla medlemsstater ?
borde inte kontrollen över verkställandet skärpas ?
skulle det inte vara lämpligt att på kort sikt , enligt exemplet från rotterdam , börja kontrollera enligt ett poängsystem , där till exempel fartygets ålder räknas in , om det är enkelväggigt eller dubbelväggigt , om det seglar under bekvämlighetsflagg .
kort sagt , kontroll av äldre fartyg under internationell standard skall ha högre prioritet än fartyg som uppfyller alla kvalitetskrav .
erika byggdes av ett japanskt skeppsvarv , enkelväggigt .
för närvarande finns ytterligare fyra systerfartyg i trafik .
bygget stoppades då för tiden på grund av att faran för rostbildning var extra stor för den typen av fartyg .
vissa av dem seglar också under maltesisk flagg .
nu väntar vi på nästa olycka .
borde det inte vidtas några sanktioner , som kommissionären sade , mot klassificeringssällskapet ?
rina har för närvarande fått dåligt rykte .
malta är på väg att inleda anslutningsförhandlingarna .
jag anser att europeiska unionen kan bevilja malta inträde endast om det finns garantier för att den maltesiska flaggan i fortsättningen kommer att segla prickfritt .
mina damer och herrar ! jag skulle uppskatta om ni ville visa litet bättre disciplin , för vi börjar bli försenade , och denna försening kommer att gå ut över den tid som är avsatt till frågestunden med frågor till kommissionen .
herr talman ! strax innan jag gick ned i kammaren fick jag ett e-mail med en ganska känsloladdad beskrivning från en svensk kvinna som hade valt att tillbringa nyårsaftonen vid den franska kusten i bretagne i stället för att vara hemma och fira med sina släktingar .
liksom många andra hundratals frivilliga hade hon sett förstörelsen , tvättat fåglar och städat upp efter de ansvariga som inte fanns vid kusten de kvällar och nätter , när de verkligen skulle ha behövts där .
som så många andra , undrar även jag var de ansvariga finns .
var finns redarna och transportbeställarna när dessa katastrofer inträffar ?
kanske vore det dags för oss att börja fundera över att inrätta en gemensam miljöbrottsmyndighet , som skulle kunna ta upp denna typ av brott .
det är inte första gången vi ser oljeutsläpp , avsiktliga eller oavsiktliga .
jag skulle vilja tacka grossetête och hennes kolleger för att de har lagt fram detta förslag för parlamentet .
brittiska massmedia har rapporterat mycket om miljökatastrofen då erika sjönk utanför bretagne och läckte ut 10 000 ton olja .
trots att storbritannien och frankrike har haft sina meningsskiljaktigheter på senaste tiden kan jag försäkra er att mitt land känner stort medlidande med alla de drabbade .
tv-bilderna av den skada er kustlinje och ert djurliv , särskilt fåglar och det redan tynande fiskbeståndet , har lidit fick oss att minnas liknande katastrofer i storbritannien , såsom torrey canyon 1967 , och har fått många britter att ställa upp med frivilligt arbete .
jag välkomnar dessa gemensamma ansträngningar att reparera skadan .
det är tydligen ett problem för hela eu : s kustlinje som kommer att kräva fantasifulla lösningar .
i stället för att låta de mest drabbade områdena och försäkringsbolag som lloyds i london bära kostnaderna för dessa katastrofer måste vi utveckla nya tekniker för att återvinna mycket mer än 10 procent av den förlorade oljan från havet .
eftersom försäkringsmarknaden betalar räkningen för närvarande finns små ekonomiska incitament för detta .
i slutändan måste den som förorenar betala .
dessutom måste vi bygga vidare på rådets direktiv om genomdrivande av internationella normer för fartygssäkerhet och förebyggande av föroreningar genom att säkerställa att målet att 25 procent av de fartyg som anlöper eu : s hamnar skall kontrolleras uppfylls och att kontrollerna håller hög standard .
dessutom anser jag , även om jag inte är emot att fartygens ägare registrerar sina fartyg i vilket land de vill , att en striktare tillämpning av internationella bestämmelser fordras .
snarare än att förbjuda bekvämlighetsflagg , vilket skulle vara ett brott mot varje suverän stats rätt att ha en handelsflotta , måste nationella sjöfartsmyndigheter i enlighet med 1995 års eg-direktiv om hamnkontroll pålägga utflaggningsländer som inte uppfyller sina åtaganden enligt internationella avtal effektivare sanktioner .
jag hoppas verkligen att kommissionen och rådet , speciellt under det franska ordförandeskapet senare i år , kommer att titta noggrant på dessa alternativ och jag rekommenderar helhjärtat parlamentet att anta denna resolution .
herr talman ! jag vill börja med att uppriktigt tacka för alla initiativ , inte bara från de olika grupperna , av grossetête och av europeiska folkpartiets grupp ( kristdemokrater ) och europademokraterna , utan även från wurtz och gruppen europeiska enade vänstern / nordisk grön vänster , till denna debatt som har gjort att vi har kunnat föra en viktig diskussion i positiv anda .
min avsikt är att lägga fram ett meddelande före utgången av mars månad , och det är möjligt att det kommer att innehålla lagtexter , det vill säga ändringar av konkreta direktiv så att en diskussion kan föras i rådet och i parlamentet .
jag skulle vilja påstå att det här i själva verket inte bara handlar om ett miljöproblem ; det är ett omfattande miljöproblem , men det är också ett omfattande socialt problem ; det finns män och kvinnor som är beroende av fångst av fisk och skaldjur , av tjänstesektorn eller turistsektorn i dessa kustområden ; det är områden som är utsatta ur miljösynpunkt , men även utsatta vad beträffar den sociala utvecklingen och den territoriella jämnvikten .
därför måste vi vara särskilt försiktiga så att vi i den mån det är möjligt undviker att en situation som denna uppstår igen .
roth-behrendt sade att ingenting har gjorts .
jag tror nog att kommissionen tidigare har gjort en del , men ännu mer måste göras .
beviset på detta är att nordamerikanerna , efter exxon valdez , inom ett år antog en lagstiftning som var extremt sträng och extremt hård , och som innebär en risk att man , som jag redan har påpekat , omdirigerar de båtar hit som inte accepteras av de nordamerikanska hamnarna .
i europa har vi , sedan amoko cadiz eller urquiola vid den spanska kusten år 1976 eller torrey canyon samma år , eller sedan alla andra fall som har förekommit , börjat lagstifta på allvar sedan år 1994 och 1995 , och i synnerhet på senare år .
de senaste åren har man dessutom poängterat säkerheten vid passagerartransporter .
enligt min uppfattning måste vi nu göra viktiga och angelägna insatser för att bemöta de nya problemen , som även härrör sig från den nordamerikanska lagstiftningen , där man poängterar säkerheten vid transport av farligt gods inom sjöfartssektorn .
mina damer och herrar , jag har tagit upp en rad frågor som vi kan gå in på mer i detalj , om ni vill , i samband med att jag infinner mig i det utskott som berörs av frågan , eller annars i samband med att jag lägger fram konkreta initiativ de närmaste månaderna .
min avsikt är - och det är något jag vidhåller - att vi påbörjar diskussionen i slutet av mars , en tidpunkt som sammanfaller med ett ministerråd , och att vi , givetvis innan det portugisiska ordförandeskapets period är till ända , får ett diskussionsunderlag .
bekvämlighetsflaggen är ett problem , men det är inte det enda .
rumänien är inte ett land med bekvämlighetsflagg , men man har ändå en mycket hög felkvot vid inspektioner . ännu högre än länderna med bekvämlighetsflagg .
malta och cypern har begärt inträde i unionen .
vi måste ställa höga krav i den här frågan och nu pågår förhandlingar om detta .
det kommer att leda till att vi får ompröva europeiska unionens register och ta upp det välkända problemet , som säkert kommer att dyka upp igen , vilket syftet är med ett gemenskapsregister .
även om jag tror att det skulle vara svårt , bör man utföra en granskning av de register som finns i europeiska unionens länder .
vad beträffar kontrollerna , så är själva kärnfrågan , det vill säga det första man måste ta reda på , hur den lagstiftning som vi förfogar över har fungerat , precis som hatzidakis påpekade .
vi har ju redan en lagstiftning .
enligt den information som kommissionens tjänsteenheter tillhandahållit mig har lagstiftningen i många medlemsstater inte tillämpats i tillräcklig utsträckning , på grund av brist på personal , resurser och inspektörer .
problemet är inte att endast 25 procent kontrolleras , utan snarare hur urvalet går till , hur man hittar de fartyg som utgör den största risken , utifrån fartygens ålder eller utifrån flaggens tidigare riskfaktor .
tyvärr gömmer sig dessa 25 procent bakom flagg som de vet kommer att uppfylla kraven : inspektionerna går då snabbare och arbetet är lättare att utföra .
därför måste man , förutom att vidta förändringar , även vidta åtgärder för att undersöka vad som redan görs , förutom några tilläggskrav beträffande granskningarna , i synnerhet i förhållande till de olika fartygens ålder .
där finns solas ( internationell konvention om säkerhet för människoliv till sjöss ) och marpol ( en internationell konvention om förhindrande av havsföroreningar från fartyg ) , två avtal inom ramen för internationella sjöfartsinspektionen , som bör göras obligatoriska i unionens samtliga stater så att man sedan kan kontrollera hur de tillämpas .
vad beträffar unionens inspektörer , anser jag att subsidaritetsprincipen motiverar att man godkänner att medlemsstaterna utför dessa inspektioner , vilket inte hindrar att kommissionen kontrollerar att staterna utför sin uppgift på rätt sätt .
slutligen vill jag poängtera ansvarsfrågan .
inte bara beträffande maxbeloppen som jag anser bör vara jämförbara med de nordamerikanska .
vi har fastställt 180 miljoner dollar ; i förenta staterna talar man om 1 000 miljoner dollar som ett tak för skadeersättning .
jag anser att vi bör höja det aktuella beloppet , så att vi närmar oss de nivåer som finns i förenta staterna , men att vi även bör kräva en omprövning av totalsumman för försäkringarna av fartygen , och därmed rederiernas ansvar , och låta ansvaret även omfatta dem som chartrar fartygen , ägarna av lasten .
så länge man inte utkräver något ansvar av de som äger lasten , mina damer och herrar , så kommer dessa problem enligt mig inte att kunna lösas .
det var allt , jag skall inte breda ut mig mer än såhär .
vi kommer att få andra tillfällen att diskutera detta .
men det är utan tvekan så att vi , som någon talare sade - och jag tackar för era inlägg som alla varit positiva och relevanta - måste förhindra att vi inom ett , två eller tre år åter står här och säger att vi inte har gjort det vi bör .
för min del kan jag , efter att ha diskuterat det med de övriga kommissionärerna , säga att kommissionen är beredd att inför parlamentet och rådet lägga fram de lagstiftningsåtgärder , ändringar och direktiv som krävs för att tillförsäkra oss den högsta möjliga säkerhetsnivån .
detta förutsätter en politisk vilja från parlamentet- och jag ser att jag kan räkna med den - liksom även från ministerrådet .
vi har med glädje noterat er samarbetsvilja .
jag har fått 8 resolutionsförslag i enlighet med punkt 2 i artikel 37 i arbetsordningen till följd av kommissionens uttalande .
stormar i europa
nästa punkt på föredragningslistan är kommissionens uttalande om stormarna i europa .
jag överlämnar ordet till barnier som företrädare för kommissionen .
herr kommissionär ! jag vill tacka för era uttalanden , särskilt de konkreta förslagen angående de olycksdrabbade som väntar sig oerhört mycket av europeiska unionen , och av det stöd som vi kan ge dem .
några dagar efter de hemska stormarna sände jag personligen en skrivelse till er , för att be er att försöka få den franska regeringen att justera mål 2-områdena , så att alla drabbade områden kan få mål 2-stöd , såväl i frankrike som i andra länder .
jag antar att det är gjort , eftersom ni inte talade om det .
vi vet att man har alla svårigheter i världen att få stöd om man inte ingår i ett mål 2-område .
det är således bättre att genast lösa det här problemet .
ni vet också att det inte endast är ett kortsiktigt problem , utan även ett problem på medellång och lång sikt .
jag skall förklara mig .
jag var i lorraine när de förfärliga stormarna skövlade omkring 20 procent av lövskogarna .
för vissa s.k. skogskommuner är skador på 20 procent en enorm förlust .
vi vet till exempel att det krävs mellan 150 och 200 år innan ett träd uppnår mogen ålder . den förlust som drabbar dessa kommuner sträcker sig således inte endast över ett , två eller fem år , utan en mycket längre period .
de berörda kommunerna uppskattar att det rör sig om 40 år .
jag anser följaktligen att det kommer att bli mycket svårt att med hjälp av bidrag kompensera dessa landsbygdskommuners intäktsförluster .
den aspekten tror jag att vi måste bära med oss och inte glömma den när vi vidtar olika politiska åtgärder .
det stämmer att skogssektorns problem är oerhört sammansatt .
ni talade om att frigöra medel för virkeslagren , eftersom priset inte får sjunka .
å andra sidan kommer även de kommuner som inte berördes av stormarna att lida skada , eftersom office national des forêts ( ung . skogsvårdsmyndigheten ) har beslutat att frysa skogsavverkningen under fyra års tid .
de kommuner som inte har lidit förluster kommer således ändå att få se sina inkomster minska .
detta säger jag för att visa er att problemet är ytterst invecklat , och jag vill än en gång tacka kommissionen för att den analyserar situationen så grundligt som möjligt .
jag skulle också vilja uppmärksamma er på det faktum att det visserligen har inträffat en ekonomisk katastrof , men att de verkliga miljökatastroferna ännu inte har inträffat .
det sade ni själv , herr kommissionär - stormarna är inte alltid naturkatastrofer , och vår bedömning är att de är ett första tecken på klimatförändringar .
vi bör därför se över vår politik för att integrera denna omständighet .
herr talman ! alla de som kom hit med bil , tåg eller flyg , har kunnat konstatera vidden av de skador som framför allt drabbat frankrike till följd av orkanen , en orkan av en aldrig tidigare skådad styrka , som slog till mot europa i slutet av förra månaden .
vad kan europaparlamentets ledamöter göra inför en katastrof av den omfattningen ?
först och främst vill jag hedra alla mina kolleger , borgmästare och förtroendevalda , som varje dag har fått lugna människor , organisera solidaritetsarbetet och samarbeta med de offentliga tjänsteföretagen .
de har gjort sig väl förtjänta av sina medborgares förtroende .
jag vill också tacka medlemsstaternas räddningstjänster och väpnade styrkor , som inom ramen för ett exemplariskt mellanstatligt samarbete kom för att stödja sina franska kollegers ansträngningar .
jag skulle också vilja fundera över den paradoxala situation vi befinner oss i när det gäller katastrofstöd .
hade denna katastrof ägt rum i guatemala eller turkiet hade vi genast kunnat ta gemenskapens budget i anspråk för att hjälpa offren , men i våra länder är inget sådant möjligt eftersom det saknas lämpliga budgetposter .
vi måste också be kommissionen att inte hindra lokala myndigheter och staterna från att bistå de företag som har drabbats av katastrofen , dvs. att inte tillämpa gemenskapens konkurrensregler på ett alltför strikt sätt .
jag tänker särskilt på de hårt drabbade fiskarna och mussel- och ostronodlarna .
som ni sade herr kommissionär , måste de få ersättning för det påtvingade verksamhetsavbrottet , och de investeringar som måste byggas upp på nytt skall kunna få stöd genom det finansiella instrumentet för utveckling av fisket ( ifop ) .
vidare tror jag inte att en automatisk tillämpning av de fleråriga utvecklingsprogrammen ( fuf ) är på sin plats i olycksdrabbade kustområden .
jag uppmanar därför kommissionen att avstå från det , för att i stället hjälpa dem som får sin försörjning av havet att göra de investeringar som nu är nödvändiga .
herr talman , kära kolleger ! de stormar som härjade i frankrike natten mellan den 26 och 27 december har som tidigare nämnts orsakat 90 döda och åsamkat skador för 75 miljarder franc , dvs. 11 miljarder euro .
knappt tre veckor efter olyckan var tusentals människor fortfarande utan elektricitet och telefon , 500 000 hektar skogsområden och 100 miljoner kubikmeter träd hade förstörts och det historiska arvet hade också skadats , vilket det sorgliga exemplet versailles slottspark vittnar om .
inför en sådan katastrof förefaller det därför naturligt att den nationella och europeiska solidariteten kommer de olycksdrabbade och de mest berörda personerna till del .
men i likhet med vad föregående talare har sagt , och vad ni , herr kommissionär , svarade min kollega jean-claude martinez angående en annan tragedi - nämligen översvämningarna i sydvästra frankrike i november månad - är det visserligen så att ni ser med oro på katastroferna , men det enda ni gör är att erinra om att budgetposten för hjälp vid naturkatastrofer har avvecklats .
detta leder oss fram till en chockerande paradox , som framhölls av föregående talare , nämligen att det är lättare , mycket lättare , att hjälpa offren för naturkatastrofer utanför unionen än på unionens territorium .
herr kommissionär ! ni begränsar er till , och vi förstår er , att erbjuda oss den hypotetiska och avlägsna möjligheten att få strukturstöd enligt det nya mål 2 eller övergångssystemet för mål 2 och mål 5b .
det var de ordalag ni använde i det skriftliga svaret till min kollega den 11 januari 2000 .
jag har en kopia till ert förfogande .
vi förstod mycket väl att ni inte kunde säga annat - inför den oansvariga attityd som inte endast är kommissionens utan också parlamentets - och att ni ingenting kan göra i brist på rättsliga och finansiella grunder .
men för guds skull , jag ber er , och det säger jag utan någon som helst ilska gentemot er , presentera inte redan tidigare planerade stöd som hjälp till stormarnas offer , de är ju stöd som går inom ramen för en regionalpolitik som inte har någonting med detta att göra .
inom ramen för en tilläggsbudget krävs det således att vi snarast återupprättar den budgetpost vi tilldelades för naturkatastrofer .
vi måste utnyttja stödmedlen från toppmötet i berlin , och vi måste ändra på den skogspolitik som bedrivs i de flesta av unionens länder , men det är ett annat problem .
herr talman , herr kommissionär , mina kära kolleger ! europa har vid detta millennieskifte utsatts för en hård prövning .
först av allt vill jag uttrycka min djupa sympati med de familjer som försänkts i sorg av de oväder som härjade i europa i december .
stormarna är en miljökatastrof utan tidigare motsvarigheter för våra skogar .
tillåt mig sända en särskild tanke till skogarna i min region , lorraine , där skadorna var avsevärda .
och jag vill gratulera de regionala myndigheterna , alla frivilliga och de offentliga företagen till deras exemplariska mobilisering . men tyvärr har de ännu inte sett ljuset i slutet av tunneln .
det är europas skyldighet att stödja dem och på så sätt komplettera de berörda medlemsregeringarnas insatser .
jag välkomnar med nöje barniers uttalande , liksom de åtgärder som kommissionen har aviserat .
jag skall inte förbigå den ekonomiska dimensionen av frågan ; skogssektorn är ödelagd och en hel befolkning lider av de tragiska konsekvenserna .
gemenskapens åtgärdsprogram för civilt skydd , vilket inrättades genom rådets beslut av den 9 december förra året , inleddes den 1 januari 2000 .
jag vill be staterna att gripa tag i det tillfället : detta program måste fungera fullt ut .
det har varit effektivt på vissa områden - och jag betvivlar inte att kommissionär barniers uttalanden är ärliga - men jag beklagar att programmen för skogsbruket fortfarande ligger i sin linda .
i väntan på att medel frigörs på gemenskapsnivå , bör man prioritera ett materiellt stöd inom ramen för medlemsstaternas partnerskap .
det är således brådskande att stärka skogssektorn och upprusta det så fort som möjligt .
lån av skogsutrustning och tillhandahållande av behörig personal ingår också i ett sådant arrangemang .
en kommande utmaning blir att undvika växtskyddsproblem som hänger samman med att stora mängder trä överges i skogen , och att grundvattnet förorenas till följd av att det skapas lika betydande virkeslager .
till sist är det absolut nödvändigt att bromsa utnyttjandet av avverkningsklara träd , och i stället främja köp av stormfällda träd .
denna virkesförsäljning bör understödjas av en omfattande medial bevakning på medlemsstatsnivå .
biståndet till uppsamling av trä utgör självklart bara ett första steg när det gäller att stödja återställandet av skogarna och den fysiska planeringen för landsbygden .
jag uppmanar kommissionen att integrera detta i ett reflektionsarbete om förvaltningen av problemen efter katastrofen .
det här är således ett sorgligt tillfälle för europa att gripa tag i , så att dess skogrikedomar förnyas och skogarna därmed kan uppfylla sin uppgift att bevara vilda djur och växter och naturliga livsmiljöer samt sin roll i våra länders ekonomi .
för stunden krävs det således en solidaritet och ett samarbete mellan medlemsstaterna inför en ekonomisk och miljömässig katastrof .
det är europas sak att föreslå prioriterade åtgärder för att rädda skogssektorn , så att denna solidaritet verkligen blir meningsfull .
orkanen &quot; lothar &quot; måste ge oss anledning att överge vår princip att uteslutande återställa det som skadats , vilket också här diskuteras i främsta hand , och i stället tillämpa försiktighetsprincipen , där även de eventuella upphovsmännen skall ställas till ansvar .
de aktuella programmen måste påskyndas .
åtagandet från kyoto kan exempelvis inte genomföras med kommissionens nuvarande koncept .
handeln med utsläppsrätter är enligt min åsikt omoralisk och löser inte problemet , utan skjuter bara upp det .
hela skattesystemet måste på medellång sikt göras ekologiskt .
genomförandet av uppgifterna i vitboken som rör förnybara energikällor , som skulle föra med sig en massiv minskning av växthusgaserna , måste påskyndas .
allt som den nya kommissionen hittills har lagt fram i denna riktning , är inte på långt när tillräckligt , utan alltför litet !
herr kommissionär , herr talman , mina damer och herrar ! hittills har lothar varit ett helt vanligt namn .
men tyvärr har lothar erhållit en beklaglig ryktbarhet .
orkanen med samma namn svepte fram över europa och krävde , framför allt i frankrike och i tyskland , men också i schweiz , talrika offer , och efterlämnade en rågata med förödelse .
vinden besegrade elmaster , tak , vägmärken och till slut också skogen .
det rör sig ju bara om uppskattningar när vi nu hör att på kort tid ca . 120 miljoner fastkubikmeter träd fällts av stormen .
jag har lyssnat mycket uppmärksamt på er , herr kommissionär , och jag välkomnar det också utomordentligt att ni kommer att ta en titt på katastrofen lokalt i frankrike och tyskland .
om schreyer nu under de kommande dagarna är i schwarzwald , kommer den enskilde jordbrukaren eventuellt att fråga hur kommissionen nu skall kunna hjälpa honom . hur skall europa kunna hjälpa mig ?
vad säger ni då till skogsägaren , när hans skog eventuellt inte ligger i mål-2-området , om hans skog inte ligger inom 5b-området ?
hur svarar kommissionen vid besöket på plats , när ni säger till skogsägaren att vi stöder vägbyggnad och dammar , vi vill bygga upp det kulturella arvet igen , vi vill komma med erbjudanden till turisterna etc ?
att detta är välmenta råd .
men jag kommer själv från en skogsfastighet i norra tyskland , och jag kan tala om att vi i vår region redan nu märker dessa enorma skador .
man fortsätter inte med den nödvändiga gallringen av skogen , skogarna sköts inte tillräckligt .
vad vi ur kommissionens synpunkt absolut behöver , är också ett ja till de nationella stöden , så att vi inte senare åter talar om några konkurrenssituationer .
herr talman , herr kommissionär , kära kolleger ! tillåt mig att till att börja med visa på två fakta .
för det första : i början av 1999 jämnade nato i frihetens namn kosovo med marken med hjälp av bomber , med deltagande av de flesta medlemsstaterna i europeiska unionen .
nu försöker vi med gigantiska insatser åter få landet på fötter och hjälpa människorna där . detta med all rätt .
för det andra : i slutet av 1999 rasade oerhörda stormar och förde med sig död och förintelse över många landsändar inom eu .
ropet på hjälp från de drabbade besvarades av kommissionen i bryssel med en axelryckning .
vi har inga medel och inga möjligheter , hette det .
detta är fel ! ingen kan heller förstå det .
och absolut inte den som känner sin existens hotad .
människorna i europeiska unionen förväntar sig solidaritet , även inom denna gemenskap .
jag säger att de har rätt till solidaritet .
europaparlamentet måste i nödens stund se till att de också får det .
jag begär av kommissionen att den inte skall vara nödbedd utan gå offren för ovädret till mötes .
kommissionen känner bättre till medel och vägar för hjälpen än alla lokala organisationer eller myndigheter .
jag ber , kära kolleger , om ert stöd för att göra klart för kommissionen att det inte så mycket är möjligheterna att hjälpa som saknas , utan den goda viljan i många ämbetsrum i bryssel !
tillåt mig ytterligare ett påpekande : när det gäller stormens följder framgår detta mindre tydligt , men olyckan med tankfartyget utanför den franska kusten gör det helt klart att vi också i en annan fråga måste hjälpa kommissionen på traven .
vi behöver inom europeiska unionen snarast få regler beträffande miljöansvar .
det går inte längre an att allmänheten får stå för de skador , som enskilda individer ofta orsakar med sina brottsliga förehavanden .
vi måste göra upphovsmännen ansvariga för alla slags skador på vår miljö .
då kommer exempelvis alla att överväga om de skall transportera olja i ett tankfartyg , som är på väg att brytas sönder .
när jag 1994 , för mer än fem år sedan , kom med i parlamentets utskottet för rättsliga frågor och den inre marknaden , fick jag ta över uppgiften som föredragande för området med miljöansvar .
sedan dess väntar jag på ett initiativ från kommissionen , som också ger mig arbete .
det är en skandal , som snabbt måste få ett slut , och jag hoppas att detta ärende inte skjuts upp än en gång i februari !
herr talman , herr kommissionär ! denna storm vid millennieskiftet bör få oss att tänka över problemen i grunden .
det står klart att människan fortfarande inte är i stånd att undvika naturkatastrofer .
det har alltid funnits och kommer alltid att finnas naturkatastrofer .
naturligtvis behövs det solidaritet i detta sammanhang .
det behövs säkerligen ett civilskydd över hela europa , och det måste också inrättas en budgetpost för naturkatastrofer i eu : s budget .
men - och det är det viktigaste - misstagen när det gäller förhållandet mellan natur och människa begås alltid av människan - även om de ofta görs över hundratals år - och aldrig av naturen , ty naturen kan inte göra några misstag .
skadorna i detta sammanhang berodde på befolkningstätheten , på infrastrukturens utformning och i fråga om skogen naturligtvis också på de många monokulturerna .
givetvis är jag positiv till att vi skall hjälpa så långt det är möjligt .
men vid hjälpen skall man beakta att el- och telenät kanske i framtiden i större utsträckning bör läggas under jord .
vi måste se till att vi får mindre kretslopp , och vid nyplanteringen av skog framför allt satsa på stabila blandskogar , och inte på monokulturer .
den viktigaste diskussionen i detta sammanhang är emellertid klimatet .
vi har hittills varit priviligierade i europa , eftersom vi har golfströmmen , och golfströmmen fortfarande fungerar .
amerika och sydostasien har det mycket sämre ställt , vad gäller klimatet och stormarna .
vi har lyckligtvis golfströmmen .
men vi lider liksom de andra också av växthuseffekten .
den har - hur svårt det än är att demonstrera klimatförändringen med hjälp av räkneexempel - delvis åstadkommits av människorna .
vi måste i större utsträckning iaktta direktiven från miljökonferensen i kyoto .
vi måste minska på koldioxidutsläppen , börja använda förnybara energikällor och i detta sammanhang generellt fråga oss , hur europas skogar mår .
herr talman ! jag anser att det i första hand är offren vi bör beklaga .
förlusterna är oersättliga .
för det andra välkomnar vi solidariteten de franska provinserna och medborgarna emellan , och övriga länders solidaritet med frankrike som är det land som har drabbats hårdast .
eftersom jag inte har så lång tid på mig , herr talman , vill jag endast ta upp två aspekter i vår resolution .
den första tycker jag att kommissionären indirekt erkänner i sitt anförande , när han ställer sig frågan om det rör sig om naturkatastrofer eller ej .
experterna blir ju ständigt mer övertygade om att det finns ett samband mellan klimatförändringarna och människornas agerande i allmänhet och det ökade antalet naturkatastrofer på senare år .
de senaste tio åren har temperaturen stigit mer än den hade gjort under den resterande delen av århundradet .
därför bör europa tydligt ta ställning för kyotoprotokollet och komma med konkreta förslag .
den andra aspekten är att det var jag som var föredragande för civilförsvaret i europa , och jag är helt enig i kommissionärens förslag att upprätta en europeisk civilförsvarsmakt .
dessutom bör man använda sig av en budgetpost utöver de vanliga , precis som en katastrofsituation är något utöver det vanliga .
först av allt skulle vi vilja uttrycka vår medkänsla med alla de familjer och samhällen som har förlorat medlemmar i denna fruktansvärda tragedi .
det är faktiskt förlusten av liv som gör denna speciella katastrof extraordinär med europeiska mått .
det är beklagligt att vi inte har några verktyg för att ge bistånd i sådana här situationer .
jag vill tacka kommissionären för hans innehållsrika uttalande i frågan och hans förslag att vi faktiskt skulle kunna organisera oss på europeisk nivå för att ge bistånd till medlemsstater och regioner som upplever liknande tragedier .
en andra sak vi bör komma ihåg är att vi hade en budgetpost tidigare .
den var mycket liten .
den räckte inte till mycket men den missbrukades flera gånger av ledamöter av denna kammare som föreslog åtgärder när katastroferna inte ens var stora .
medlemsstaternas tjänstemän och ministrar kom till bryssel , viskade med kommissionen , fick några euro och en politisk poäng genom att de hemförde stöd till sina valkretsar .
så det var inte många som sörjde att denna budgetpost avskaffades .
jag tror att vi bör återinföra denna budgetpost .
när vi hade jordbävningen i grekland , som var en stor katastrof , hade inte gemenskapen något instrument för att visa grekerna sitt medlidande och sin solidaritet .
detsamma gällde när översvämningarna drabbade frankrike , och detsamma händer nu igen .
dessa katastrofer är stora , vi borde ha ett instrument men vi har det inte .
vi bör återinföra detta instrument och göra reglerna strikta , så att vi bara använder detta speciella instrument i situationer då allvarliga katastrofer inträffar .
vi kan spara det från år till år och tillse att vi har ett instrument för att handskas med stora olyckor när de inträffar .
i irland var det inte så illa den här gången , även om vi har haft många allvarliga stormar på atlanten .
vi hade översvämningar i irland också och jag vill ge uttryck för min medkänsla med de människor i irland som drabbades av dessa .
mina kära kolleger ! det får inte bli så att var och varannan bland oss tappar minnet .
det stämmer att kommissionen och parlamentet fattade ett gemensamt beslut , vilket syftade till att avskaffa budgetposterna för katastrofhjälp .
det stämmer att det finns mycket europeiska pengar - kommissionär barnier har pekat på att han kommer att utnyttja artikel 30 i arbetsordningen om landsbygdens utveckling för ostronodlingarna och jordbruket ; artikel 33 för skogsbruket ; undantagen till konkurrensreglerna i artikel 87.2 i fördraget för företagens del samt strukturfonderna för offentliga anläggningar .
ändå kvarstår det faktum att det i dag inte uppbringas ett enda öre mer än vad som skulle ha tilldelats före stormen , för att uttrycka en konkret och aktiv solidaritet .
för staterna gäller det helt enkelt att agera kommunicerande kärl och ta från ett ställe för att ge till någonting annat .
detta är otillräckligt , och därför gläder det mig personligen att barnier tog upp den idé som ligger mig varmt om hjärtat , en idé jag för övrigt framförde när jag uttryckte mina önskningar till pressen i bordeaux , nämligen inrättandet av en förstärkt politik för ett europeiskt civilskydd .
jag tror att medborgarna måste uppleva våra omedelbara åtgärder som påtagliga , om vi vill att det för oss så eftersträvansvärda europeiska medborgarskapet skall existera , och om vi vill att det mandat som vår talman fontaine har ställt upp skall bli verklighet , dvs. att unionen och europas medborgare skall närma sig varandra .
jag tror därför att en europeisk civil säkerhetsstyrka borde vara något för oss att sträva efter ; att vi upprättar en formering av blå baskrar för civil säkerhet som skall vara närvarande på platser med svårigheter - inom unionen för att vi i dag inte har någon katastrofstrategi , men vid behov också utanför unionen , till exempel i venezuela eller andra länder .
jag vill också säga kommissionär barnier att han i mig har en allierad som agerar för den här idén , som jag anser vara generös och europeisk .
herr talman , herr kommissionär , kära kolleger ! jämfört med hur ofta det uppträder stormar i andra områden i världen , är vi i europa relativt förskonade .
trots detta har stormarna under den sista decemberveckan visat vilka följder de kan få , och att vi också kommer att få stora problem .
alla som åkte till strasbourg med bil eller järnväg kunde övertyga sig om hur stormen rasat också i alsace .
jag vill därför uttala min medkänsla med alla medborgare i de regioner där stormen rasade så vilt , och samtidigt här i kammaren påpeka vikten av att stödja regionerna och människorna .
vi alla vet att det i morgon lika gärna kan vara en annan region i europa som drabbas på liknande sätt .
det gäller nu att så snabbt som möjligt ta till vara dessa vindfällen .
ty var och en vet att vi kan drabbas av ännu större katastrofer , om vindfällena får ligga kvar för länge i skogen .
det måste också påpekas att exempelvis barkborren finner den bästa grogrunden för sin utbredning och för sina larver i vindfällena , och att det därigenom orsakas följdskador , som vi i dag ännu inte kan få någon uppfattning om .
därför är det absolut nödvändigt att ta till vara vindfällena redan innan den varma årstiden börjar .
den verkliga omfattningen av skadorna inom skogsbruket kommer vi att få reda på först om tiotals år .
ty vi vet alla hur lång tid ett träd behöver på sig för att växa .
här räknar man i årtionden , och inte i år .
dessutom vill jag påpeka att det inom skogsbruket säkert inte bara gäller träproduktion , utan att de skyddade och de skyddande skogarna är en väsentlig faktor i vissa regioner .
jag vill därför med stolthet säga att de österrikiska utbildade skogsarbetarna också är beredda att ...
herr talman ! vår djupaste medkänsla går till alla dem som drabbades av stormarna .
ibland är vi inom gemenskapen egentligen inte medvetna om vad som händer i andra länder .
i irland var mediatäckningen av det sjunkna tankfartyget väldigt liten .
jag ombads berätta om konsekvenserna av stormarna i irland .
vi hade stark vind och ett långvarigt skyfall utan motstycke som lades till de svårigheter som redan fanns och resulterade i att hundratals hektar översvämmades och ibland lades under så mycket som 45 centimeter vatten .
vi upplevde den mänskliga misären med översvämmade hem och gårdar , utan hälsovård och dricksvatten , och de miljömässiga katastroferna med e-kolibakteriesmittat vatten .
jag talade med jordbrukare vars tackor fick missfall efter att ha druckit av det infekterade vattnet .
naturliga livsmiljöer förstördes .
därför ber jag er komma ihåg irland i detta speciella fall .
jag tackar kommissionären och stöder honom mycket starkt vad gäller hans europeiska insatsstyrka .
herr talman , herr kommissionär , mina damer och herrar ! jag ansluter mig till alla dem som har uttalat sin solidaritet med offren för stormen .
jag vill också än en gång peka på betydelsen för skogsbruket i hela europa .
ty vi kommer ju att i alla områden i europa få massiva effekter på skogsbruket , och jag tror att man här långsiktigt måste överväga hur man skall hantera sådana problem i framtiden .
vi vill säkert inte ha någon organisation av marknaden för skogarna , men vi måste eventuellt skapa ett system , kanske även i samarbete med de privata försäkringsbolagen , och tillsammans med dem på något vis mildra sådana effekter för dem som drabbats .
vi kommer tyvärr även i framtiden att tvingas räkna med dylika svåra katastrofer .
det finns sådant som tyder på det , det har redan berörts här , det finns inga bevis , men tecken som tyder på att det ökande antalet stormar över hela världen har att göra med miljökastastrofen .
forskarna är naturligtvis ännu inte eniga . men de flesta är relativt säkra på att om vi fortsätter med utsläppet av växthusgaserna så kommer dessa stormar naturligtvis att drabba oss ännu hårdare i det århundrade som just har börjat .
jag tror att vi än en gång bör erinra om ett förslag som väcktes av en tidigare kollega till oss , tom spencer , här i kammaren ; enligt det bör vi inte ge stormarna några kvinnliga eller manliga förnamn , utan döpa dem efter dem som orsakar växthuseffekten - han nämnde då oljekoncernerna .
här bör man dock säkerligen undanta shell och bp , eftersom de har ändrat sin politik och inte bara satsar på försäljning av miljöskadliga fossila bränslen , utan också investerar i framtidsdugliga energiformer .
detta sammanhang måste vi inse ; jag håller inte med dem som schablonmässigt säger att växthuseffekten bär skulden för denna storm , men att vi måste befara ytterligare katastrofer , om vi inte snabbt växlar spår , det är relativt säkert !
livsmedelssäkerhet
jag har erhållit sju resolutionsförslag som lagts fram i enlighet med artikel 37.2 i arbetsordningen . nästa punkt på föredragningslistan är meddelande om livsmedelssäkerhet och uttalande av kommissionen .
herr talman ! det gläder mig mycket att kunna ta detta första tillfälle i akt att tillsammans med min kollega liikanen för parlamentet dra upp huvudlinjerna i kommissionens vitbok om livsmedelssäkerhet , som antogs i onsdags , 12 januari .
vid min utfrågning i september lovade jag att denna vitbok skulle levereras snabbt .
jag är glad att vi har kunnat leverera den så snabbt .
mellan tre och fyra månaders intensivt arbete sedan den nya kommissionen utsågs i september ligger till grund för vitboken .
den bygger på de omfattande rådslag som har förekommit under de senaste åren sedan kommissionens grönbok om livsmedelslagstiftning utkom .
den avspeglar också våra erfarenheter från nyligen aktuella larmrapporter om sådant som dioxin och slam liksom från bse-krisen .
vitboken avspeglar också detta parlaments intressen , vilka ni har beskrivit både för ordförande prodi och för mig vid de många tillfällen då vi har debatterat livsmedelssäkerhet i denna kammare sedan kommissionen utsågs .
jag behöver inte påminna er om att konsumenternas förtroende för europas livsmedelssäkerhetssystem allvarligt har påverkats av kriser och larmrapporter under de senaste åren och månaderna .
kommissionen har förbundit sig att återskapa detta förtroende genom att skapa världens mest moderna och effektiva system för livsmedelssäkerhet .
när jag lanserade vitboken förra veckan sade jag att kundvagnen är ett av de mest kraftfulla vapnen på denna jord .
europas konsumenter fattar de mest omdömesgilla besluten .
om deras förtroende rubbas avspeglar inköpsbesluten detta .
detta har i sin tur dramatiska konsekvenser för jordbrukare , producenter och industrin i allmänhet .
i en bransch som omsätter omkring 600 biljoner om året kan även en liten nedgång i förtroendet få betydande konsekvenser .
inom den agrara livsmedelssektorn och jordbrukssektorn finns över 10 miljoner anställda .
ett högt förtroende är en förutsättning för att öka sysselsättningen och konkurrenskraften .
denna förtroendekris har också fått den olyckliga men oundvikliga konsekvensen att konsumenternas förtroende för system och institutioner på nationell och europeisk nivå som skall övervaka och säkerställa högsta möjliga livsmedelssäkerhet har försvunnit .
när jag säger allt detta vill jag också slå fast att europa trots detta har en av världens bästa livsmedelsindustrier och också ett av de säkraste systemen för livsmedelskontroll .
utmaningen är att göra systemet till de allra bästa .
det övergripande syftet med vitboken om livsmedelssäkerhet är därför att skapa erforderlig lagstiftning och strukturer som kan garantera konsumenterna högsta möjliga hälsoskydd vid livsmedelskonsumtion .
vi sätter upp en krävande och ambitiös dagordning för förändring .
kommissionen kommer att behöva parlamentets fulla stöd om vi skall kunna uppnå våra mål enligt tidsplanen .
vi kommer också att behöva rådets och andra nyckelfunktioners fullaste stöd .
i vitboken om livsmedelssäkerhet beskrivs en omfattande uppsättning åtgärder som fordras för att komplettera och modernisera dagens livsmedelslagstiftning inom eu .
alla dessa åtgärder syftar till att göra den mer konsekvent , begriplig och flexibel .
vi vill verka för en bättre tillämpning av denna lagstiftning och ge konsumenterna större öppenhet .
i den detaljerade handlingsplanen om livsmedelssäkerhet i vitboken finns en preciserad tidtabell för åtgärderna under de närmaste tre åren .
över 80 åtgärder planeras .
vårt mål är att ha skapat en konsekvent och modern livsmedelslagstiftning vid utgången av år 2002 .
vi planerar också att etablera en europeisk livsmedelsmyndighet år 2002 , som ett viktigt komplement till den nya livsmedelssäkerhetslagstiftningen .
denna idé kommer att bli föremål för mycken analys och debatt .
den har redan gett upphov till många kommentarer , inklusive reaktioner från parlamentsledamöter .
det kapitel i vitboken som handlar om att skapa en europeisk livsmedelsmyndighet är klart utformat för att locka fram åsikter och kommentarer .
vi vill ha in synpunkter på våra planer före slutet av april .
jag kommer att återkomma till detta rådslag om några ögonblick .
kommissionen anser att det krävs en övergripande strukturell förändring av vårt system för livsmedelssäkerhet för att säkerställa de nära besläktade målen att garantera högsta livsmedelssäkerhet och återställa konsumenternas förtroende .
varför skulle en europeisk livsmedelsmyndighet vara en viktig del av denna förändring ?
den första nyckelfrågan är oberoende .
huvudaktörerna , däribland konsumenterna , söker ett system som är oberoende och som upplevs som fristående från alla lagstadgade intressen .
vi måste också garantera förträfflighet och öppenhet .
vi har gjort många framsteg under de år som har gått sedan det reformerade systemet med vetenskapliga råd antogs som en konsekvens av bse-krisen .
emellertid menar kommissionen att vi måste gå längre .
vi måste skapa ett permanent och verkligt oberoende , utmärkt och öppet system för riskvärdering .
myndighetens huvuduppgift kommer att vara riskvärdering inom livsmedelssäkerhetsområdet .
vi tänker oss att de uppgifter de befintliga fem vetenskapliga kommittéerna som sysslar med livsmedelssäkerhet har skall överföras till myndigheten .
de kanske inte överflyttas med sin nuvarande form eller struktur - detta är en fråga som vi vill ha synpunkter på innan vi framlägger våra slutliga förslag om att inrätta myndigheten .
om vi emellertid bara skulle föreslå en ommöblering skulle detta naturligtvis inte vara tillräckligt .
som klargörs i vitboken måste den nya myndigheten ge ett mervärde .
jag anser att det nuvarande systemet med vetenskapliga råd behöver förstärkas .
inom denna myndighet tänker jag mig ett mycket starkare vetenskapligt och annat stöd för de oberoende vetenskapsmännen .
jag förställer mig också att myndigheten kommer att vara mycket mer förebyggande än vårt nuvarande system - att förekomma snarare än reagera , att identifiera frågor innan de blir till kriser .
detta förebyggande tillvägagångssätt bör bli myndighetens ledstjärna .
för att myndigheten skall kunna förebygga identifieras i vitboken ett antal nya områden som den skulle hantera .
här ingår en omfattande informationsinsamling och övervakning , samordning av vetenskaplig information inom eu och uppbyggande av starka nätverk med livsmedelssäkerhetsenheter och -organ i medlemsstaterna .
vi tänker oss också att myndighetens befogenheter skall omfatta driften av ett utbyggt snabbvarningssystem för problem med livsmedel och foder .
kommissionen har beslutat att det varken är lämpligt eller möjligt att överlåta riskhantering till myndigheten .
vi anser att beslut som gäller riskhantering fortfarande skall förbehållas kommissionen , parlamentet och rådet .
jag ber inte om ursäkt för denna inställning för jag är övertygad om att den är riktig .
naturligtvis finns det de som skulle hävda att vi bör ge en sådan myndighet lagstiftande makt .
jag accepterar inte detta synsätt och tillbakavisar det med viss hetta .
så sent som förra året ändrades fördraget så att parlamentet fick en mycket större roll i lagstiftningsprocessen .
att i detta skede ge en myndighet denna roll vore enligt min mening ett steg tillbaka och skulle innebära en urvattning av det demokratiska ansvaret .
jag är mycket intresserad av att höra parlamentets synpunkter i denna fråga .
det finns också de som hävdar att kommissionen egentligen skulle kunna ignorera den nya myndighetens råd .
jag tillbakavisar även detta resonemang .
hur kan en kommissionär för hälsa och konsumentskydd avslå eller ignorera välgrundade vetenskapliga råd från oberoende källor om livsmedelssäkerhet ?
skulle detta ligga i europas medborgares intresse ?
enligt min åsikt skulle de flesta definitivt inte göra det , om inte ett sådant tillbakavisande av de vetenskapliga argumenten hade sunda skäl , kunde försvaras rationellt och var helt rättfärdigat .
det är svårt att tänka sig en sådan situation .
jag kan försäkra er här i dag att kommissionen kommer att ta full hänsyn till myndighetens vetenskapliga råd när den utövar sin riskhanteringsfunktion .
jag har redan sagt att myndigheten kommer att ansvara för att utveckla nätverk med nationella livsmedelssäkerhetsenheter och -organ i medlemsstaterna .
detta är en stor uppgift .
vi måste utveckla en större säkerhet i den vetenskap som bär upp livsmedelssäkerheten i europeiska unionen .
myndigheten måste bli en auktoritet för vetenskaplig rådgivning och information om livsmedelssäkerhet .
denna situation skapas inte genom myndighetens blotta tillkomst utan kommer att framträda efter hand i takt med att självförtroendet stiger inom myndigheten själv .
jag tror inte att vi kan vara föreskrivande gentemot vetenskapen och råd som grundas på vetenskap .
i och med att dynamiska nätverk utvecklas med nationella livsmedelssäkerhetsenheter och -organ kommer dock myndigheten att bli dominerande på den europeiska scenen .
jag vill också gärna höra parlamentets synpunkter på detta .
som en integrerad del i en mervärdesstruktur föreslås i vitboken att myndigheten skall ha en huvudroll inom riskkommunikation : att sprida komplicerad vetenskaplig information på ett konsumenttillvänt sätt , att vara den självklara och oundgängliga instans man vänder sig till för de allra senaste riskuppgifterna , att vara mycket synlig , att berätta goda nyheter om livsmedel , att vara förebyggande .
vitboken innehåller också mycket viktiga förslag vad kontrollen beträffar .
detta är en enormt viktig beståndsdel i systemet av avprickning och avrapportering för att tillse att medlemsstaterna och aktörerna uppfyller gemenskapens lagstiftning .
jag vill se en riktig inre marknad i funktion på kontrollområdet .
i detta sammanhang föreslår vi också att den kontrollfunktion som utövas av kontoret för livsmedels- och veterinärfrågor i dublin stärks betydligt .
denna reviderade gemenskapskonstruktion skulle ha tre grundstenar : operativa kriterier som fastslås på gemenskapsnivå , riktlinjer för gemenskapskontroll och ett ökat administrativt samarbete för att utveckla och bedriva kontroll .
som en del av våra förslag på detta område - som jag har för avsikt att lägga fram mot slutet av året - kommer jag att granska om kommissionen behöver ges ytterligare maktmedel som komplement till förfaranden vid överträdelser .
dessa skulle kunna inkludera att innehålla finansiellt stöd från gemenskapen eller att återkräva medel som redan överlämnats till en medlemsstat .
dessa förslag skall ses som en del i vår strävan att ha världens strängaste normer för livsmedelssäkerhet , öka konsumenternas förtroende och vidga marknaderna för jordbrukare och producenter i unionen .
förutom förslagen om en ny europeisk livsmedelsmyndighet och ett förstärkt kontrollsystem på gemenskapsnivå innehåller vitboken förslag till en handlingsplan med ett brett spektrum åtgärder för att förbättra gemenskapens lagstiftning och göra den mer konsekvent , vilka täcker alla aspekter av livsmedelsprodukter från bondgården till köksbordet .
här beskrivs över 80 enskilda åtgärder som planeras under den period vi har framför oss i syfte att täppa till de identifierade kryphålen i dagens lagstiftning .
den nya rättsliga ramen kommer att omfatta djurfoder , djurens hälsa och välfärd , hygien , föroreningar och residuer , nya födoämnen , tillsatser , smakämnen , förpackning och bestrålning .
den kommer att innehålla ett förslag till generell livsmedelslagstiftning som inbegriper principerna om livsmedelssäkerhet såsom fodertillverkares , jordbrukares och livsmedelshanterares ansvar , om att foder , livsmedel och ingredienser skall kunna spåras , om ordentlig riskanalys genom till exempel riskvärdering - det vill säga vetenskaplig rådgivning och informationsanalys - om riskhantering - det vill säga reglering och kontroll - riskkommunikation och tillämpning av försiktighetsprincipen om och när det är lämpligt .
vad försiktighetsprincipen beträffar kan jag tillägga att kommissionen för närvarande håller på att slutföra ett meddelande som jag förväntar mig skall antas mycket snart .
jag ser fram emot ett nyttigt utbyte av åsikter i eftermiddag med parlamentets ledamöter , som förstås skulle ha föredragit att göra detta förra veckan om något lämpligt parlamentsforum hade funnits tillgängligt .
mot bakgrund av mina kontakter med ordförandena i berörda utskott inser jag emellertid att detta inte lät sig göras .
men jag vet också att vi kommer att få många fler tillfällen att överväga förslagen om en myndighet i vitboken under de kommande månaderna .
vi har nu ett antal månader på oss för att avhålla den nödvändiga debatten om kommissionens idéer om vitboken om inrättandet av en europeisk livsmedelsmyndighet .
parlamentet kommer att spela en viktig roll i denna debatt .
parlamentet spelade en avgörande roll i europas svar på bse-krisen .
det har varit särskilt aktivt sedan dess för att sätta medborgarnas oro om livsmedelssäkerheten i förgrunden .
jag väntar mig att parlamentets bidrag till debatten om myndigheten skall bli lika betydande och konstruktivt .
även om vi har ett antal månader på oss till slutet av april för att debattera denna fråga och samla in våra synpunkter inser jag fullkomligt att detta också är en mycket stram tidtabell .
jag skulle därför vilja be parlamentet att vidta lämpliga åtgärder för att tillse att dess åsikter formuleras så snabbt som möjligt .
det är viktigt att kommissionen får dra nytta av parlamentets bidrag till formandet av det som är tänkt att bli en viktig del i arbetet för att föra upp skyddet av konsumenternas hälsa till ett nytt plan och därigenom återställa konsumenternas förtroende för europeiska unionens politik för livsmedelssäkerhet .
den europeiska livsmedelsmyndigheten kommer att bli en huvudaktör i eu : s politik för livsmedelssäkerhet under kommande år .
det är viktigt att vi ger den rätt ingredienser .
herr talman ! jag tackar kommissionären för hans uttalande .
jag skulle vilja uttrycka min uppskattning av den arbetsfördelning ni har gjort och av att livsmedelsfrågorna kommer att förbli en angelägenhet för de europeiska institutionerna , inklusive kommissionen och parlamentet .
detta är alldeles rätt inställning .
men det finns ett ord som jag inte har hört er nämna i kväll .
jag hoppas att vi kan reda ut det här .
vi behöver en livsmedelslagstiftning , som ni sade , och vi behöver komma överens om detta .
det är väldigt viktigt att vi inbegriper ansvaret i denna process .
det är detta ord jag menade .
problemet hittills är att skattebetalarna har betalat när någonting har gått fel .
när vi har en kris måste vi klart slå fast i förväg att om det finns ett problem är de som är upphov till det betalningsansvariga .
herr talman ! det var en mycket bra vitbok , det vill jag inte förneka .
mina frågor gäller positivlistan för djurfoder .
det är oklart i er vitbok .
hur ser er tidsplan ut , hur snabbt kommer ni att lägga fram en positivlista ?
när kommer det att ställas samma krav på djurfoder och uppfödning som på tillverkning av livsmedel och kontroll av livsmedelstillverkningen ?
den sista delen av min fråga : när kommer bse-tester att bli obligatoriska i alla medlemsländer ?
även där är ni , beträffande förpliktelsen , något oklar i er vitbok .
tack för ert uttalande , herr kommissionär .
jag anser att de linjer ni har dragit upp vad beträffar livsmedelssäkerhetsmyndigheten speglar verkligheten .
medlemsstaterna skulle inte acceptera ett reglerande organ , så det är ingen större idé att ni föreslår ett .
för vissa delar av livsmedelsindustrin krävs uppenbarligen bättre lagstiftning och detta står klart i fråga om livsmedel och djurfoder .
i egenskap av ordförande i ett utskott som verkar komma att ägna sig nästan uteslutande åt livsmedel under de kommande tre åren måste jag dock fråga : om europa har det säkraste systemet för kontroll av livsmedel , som ni sade , varför behöver vi då 24 nya direktiv och förordningar och 20 nya ändringsdirektiv ?
för det andra , kommer inte detta att förvärra problemet med för mycket reglering från bryssel och för litet tillämpning i medlemsstaterna ?
vi ser fram emot en givande dialog med er om detta .
vad utvidgningen beträffar : vilka planer har kommissionen på att dra in ansökarländerna i debatter om dessa nya lagar , under förutsättning att kommissionen verkligen förväntar sig att de lagar som planeras i vitboken skall utgöra en del av gemenskapens regelverk senast år 2003 ?
herr talman ! först av allt skulle jag vilja tacka ahern , roth-behrendt och jackson för deras stöd för vitboken .
det tycker jag är uppmuntrande och jag ser fram emot ytterligare diskussioner med dem och med andra parlamentsledamöter om de frågor de tog upp .
ahern tog upp frågan om ansvar .
detta tas naturligtvis inte upp särskilt i vitboken förutom hänvisningen till det faktum att vi kommer att skapa bestämmelser - och det finns redan några - om möjligheterna att spåra livsmedel .
när väl detta är gjort kan frågor som ansvar tas upp .
jag har trots min bakgrund inte helt och i detalj övervägt frågor som sammanhänger med och omger ansvarsfrågorna , men jag tror att det mycket väl kan vara subsidiaritetsfrågor involverade .
men jag har noterat ert förslag och kommer att överväga det ytterligare .
roth-behrendt frågade mig om upprättandet av en positiv lista .
det är en av de frågor vi tar upp i bilagan till lagförslaget och avsikten är att upprätta en positiv lista för fodermaterial .
för närvarande är listan , som jag säger , en negativ lista som fylls på vid behov .
upprättandet av den positiva listan är en av de frågor som behandlas i bilagan som har ett datum åsatt , år 2002 faktiskt .
det snabba varningssystemet för foder är någonting vi har identifierat som en lucka i lagstiftningen .
snabb varning finns för livsmedel men inte för foder .
detta är olyckligt och det är fel , och vi tror att det är viktigt att påpeka det och införa lagstiftning som täpper till denna lucka , och detta skall göras .
medlemsstaternas arbete med bse och införandet av stickprovstest för att identifiera infektionsnivåer i medlemsstaterna pågår . jag vet att roth-behrendt har frågat mig om detta förut och jag sade att jag tyckte att det gick snabbt framåt , men jag har förstått att ärendet befinner sig på intern remiss i kommissionen och att arbete pågår .
jag hoppas att jag nästa gång ni ställer frågan kommer att vara i stånd att ge er mer detaljerad information .
jackson inriktade sig på det faktum att det finns 24 nya och 20 ändringsakter i lagstiftningen och frågar om detta innebär överreglering .
jag skulle vilja säga att de rättsakter vi har skiljt ut syftar till att täppa till luckor i gällande lagstiftning .
det handlar inte så mycket om att skapa nya system för ytterligare reglering , även om detta är en del av det , utan om att identifiera var det finns luckor och kryphål i kedjan från bondgård till middagsbord och täppa till dem .
det finns en hänvisning till ansökarländerna och detta är någonting vi tänker på .
normer för livsmedelssäkerhet och också andra säkerhetsfrågor är naturligtvis av avgörande betydelse för utvidgningen och detta är en fråga jag har tagit upp med verheugen .
herr kommissionär ! vissa medlemsländers okunnighet har fört oss in i en stor livsmedelskris i europa , och jag är , tyvärr , än en gång irriterad över att rådet i sin helhet återigen saknas i dag , när ni lägger fram detta intressanta meddelande .
jag skulle gärna vilja höra av er hur ni skall se till att en sådan ny myndighet , vad den än må heta i detalj , även får inflytande på rådet , vem i denna myndighet som skall bestämma , och vem som skall dela ut uppdragen .
naturligtvis får vi inte föreskriva något om innehållet , men jag insisterar redan på att parlamentet efter maastricht och amsterdam skall behålla sin rätt och rent av bygga ut den .
jag är mycket oroad över att vi återigen kan få en myndighet , som flyger anonym som en satellit över europa ; en sådan myndighet skulle jag älska lika mycket som djävulen älskar vigvattnet . jag hoppas att det inte kommer att ske !
även jag välkomnar vitboken .
men planerar ni att livsmedelssäkerhetsmyndigheten skall ha tillräcklig makt för att förhindra något liknande det köttkrig vi har haft och frankrikes vägran att häva importförbudet ?
ni nämnde att kommissionen har möjlighet att hålla inne anslag och bidrag för länder som agerar på det sätt som frankrike agerar .
skulle ni då också föreslå att kommissionen kan göra interimsbetalningar till exempel , liknande de brittiska jordbrukare ber om för närvarande ?
herr talman , herr kommissionär ! vid ett informationsmöte i förra veckan sade ni att eu : s livsmedelsmyndighet enligt er uppfattning inte borde förläggas på en avlägsen ort , men ni sade inte vad ni menade med denna avlägsna ort .
den verksamhet som eu-enheten i dublin bedriver har exempelvis visat att det geografiska avståndet i dag inte är något hinder för effektiv påverkan och kontakt .
man har sagt att den kommande livsmedelsmyndighetens viktigaste uppgifter är att samla in , publicera och samordna data , utfärda rekommendationer i syfte att utveckla livsmedelssäkerheten och - som ni konstaterade - samla in vetenskapliga yttranden och göra informationen lättillgänglig och lättförståelig för konsumenterna .
allt detta kan med hjälp av dagens teknik skötas var som helst inom europeiska unionens område .
jag frågar därför , vad grundar ni er uppfattning om lokaliseringen på ?
. ( en ) vad beträffar myndighetens utformning : för det första kommer den att anställa egna vetenskapsmän som kommer att hålla kontakt med och rådfråga vetenskapsmän som är experter på de just de områden som för tillfället är aktuella .
dessutom kommer livsmedelssäkerhetsmyndigheten att ha en styrelse .
ni kommer att märka av vitboken att vi inte har gått in på detaljer om hur denna styrelse skall vara sammansatt .
detta är en fråga som jag förväntar mig att parlamentet och kommissionen kommer att diskutera under de kommande veckorna och månaderna .
jag föreställer mig att styrelsen kommer att bestå av finansiärerna eller av företrädare för dessa .
i det förslag jag skall lämna till kommissionen i september måste dess funktion beskrivas i detalj .
vi har inte gjort det än , men det kommer att göras i september .
jag väntar mig inte att styrelsen skall tala om för vetenskapsmännen hur de skall sköta sitt arbete .
det skulle eliminera de vetenskapliga rådens oberoende .
men den kommer att ha en generell befogenhet , särskilt till exempel för att kräva att myndigheten granskar vissa områden som behöver utforskas .
florenz frågar om parlamentet kommer att ha någonting att säga till om här .
det är en fråga att överväga och diskutera .
det kan finnas ett antal åsikter om det .
vissa kanske intar ståndpunkten att det vore olämpligt att parlamentet eller parlamentsledamöterna - eller rent av av parlamentet utsedda ledamöter - sitter med i styrelsen .
andra kanske anser att det skulle vara en nyttig övning om parlamentet , via ombud eller ledamöterna själva , skulle få en möjlighet att diskutera vilka frågor som skall undersökas .
det tål att tänka på , men det är inte uteslutet .
florenz tog också upp frågan om anonymitet .
jag är glad att han tog upp den eftersom det är särskilt viktigt att denna myndighet har en hög profil .
den måste synas .
den måste vara känd .
konsumenterna i europeiska unionen måste veta att livsmedelsmyndigheten finns .
myndighetens vd bör vara någon som är känd , någon som kanske regelbundet medverkar i tv-program om livsmedelsfrågor , särskilt vad gäller de goda livsmedelsnyheterna om näringsvärden , kosthållning och liknande , så att konsumenterna känner till att en sådan myndighet finns om en ny livsmedelskris uppstår .
de skall vara medvetna om att de har hört talas om myndigheten tidigare under andra omständigheter och förhoppningsvis ha ett grundförtroende som redan har byggts upp genom myndighetens uttalanden .
det är därför av avgörande betydelse att myndigheten inte är anonym .
jag kommer att göra allt som står i min makt för att verka för att myndigheten får denna höga profil .
lynne frågar om myndigheten kommer att ha tillräcklig makt .
jag misstänker att frågan gäller var myndighetens befogenheter börjar och slutar och var livsmedelssäkerhetsmyndigheter i medlemsstaters ansvar och behörighet börjar och slutar .
det skulle krävas en växelverkan på vetenskaplig nivå .
det vore helt klart inte önskvärt med en situation där det uppstår motsättningar mellan vetenskapsmän som arbetar för eller är konsulter till livsmedelssäkerhetsmyndigheten på gemenskapsnivå och någon vetenskaplig åsikt på medlemsstatsnivå .
detta är en icke önskvärd situation , en situation vi inte vill se i framtiden .
det finns ett antal saker som undergräver konsumenternas förtroende , och informationsbrist är en av dem .
men information som innehåller grundläggande meningsskiljaktigheter mellan vetenskapsmän i viktiga frågor som gäller livsmedelssäkerhet är också något som inger stor oro .
vi måste försöka undvika detta och skapa strukturer som säkerställer att det finns ett ordentligt informationsutbyte mellan vetenskapsmännen , att rådslag och diskussioner genomförs till fullo och att myndigheten på gemenskapsnivå har möjlighet och mandat att fråga oberoende vetenskapsmän i alla medlemsstaterna och kanske rent av längre bort , när experter finns annorstädes , om råd och åsikter .
med tiden kommer , som jag sade nyss , inte bara myndigheten att få en tydligare profil utan dess expertis , dess moraliska auktoritet , kommer att öka i takt med att tiden går så att dess åsikter accepteras och inte ifrågasätts .
denna situation kan vi uppnå med tiden .
man kan inte lagstifta fram konsumenternas förtroende .
det är någonting man vinner med åren .
kommissionen kommer emellertid att ha möjlighet att tillse att myndighetens åsikter i vetenskapliga frågor genomdrivs genom att lagstiftning antas , vilket är kommissionens , parlamentets och rådets funktion .
jag inser att detta är en något tidsödande övning , men trots detta anser jag att införandet av lagstiftning som härrör ur myndighetens ståndpunkter är rätt väg att gå .
om lagstiftningen inte följs kan detta hanteras i domstolarna på normalt sätt .
en av de frågor som vi kan komma att tvingas ta upp med tiden är frågan om svarstider under sådana omständigheter .
jag tänkte se om någonting kan göras , så att vi får snabbare respons från domstolsprocessen .
vad gäller anslag och bidrag : ja , vi har tagit hänsyn till denna fråga .
den kommer att kräva juridisk rådgivning och detta kommer vi att begära , särskilt med tanke på att det kan ge ett snabbt svar på underlåtenhet att uppfylla gemenskapslag i avvaktan på ett domstolsutslag .
vad gäller lynnes fråga om interimsbetalningar : detta är en fråga som mycket väl kan tas upp i parlamentet , eftersom den gäller budgetfrågor .
myller frågade sedan om myndighetens placering .
inget beslut har fattats om detta annat än att säga att det är mer troligt att myndigheten placeras centralt än perifert .
jag inser att feo är placerat i dublin och , trots att jag själv kommer från den delen av världen , måste jag acceptera att det inte är europas centrum !
men feo befinner sig i en helt annan situation än livsmedelssäkerhetsmyndigheten .
feo består av oberoende vetenskapsmän och veterinärer och så vidare som reser från någon plats där det finns en flygplats - och det har vi helt klart i dublin .
livsmedelssäkerhetsmyndigheten har en helt annan situation .
den måste finnas nära kommissionen till följd av behovet av samverkan mellan de vetenskapsmän som arbetar för livsmedelssäkerhetsmyndigheten och de av oss som är involverade i lagstiftningsinitiativ .
en viktig del av kommunikationen mellan de två institutionerna kommer självfallet att bli att tillse att de av oss som sysslar med att göra upp lagförslag tydligt och klart förstår vad vetenskapsmännen menar , vilka problem de har identifierat , vilken lagstiftning som krävs för att ta itu med de frågor de tar upp .
på samma sätt kommer vetenskapsmännen att vilja ha något inflytande på utformningen av politik och lagstiftning för att tillse att lagstiftningen botar det onda de har identifierat .
jag tycker det verkar önskvärt att en sådan myndighet är centralt placerad .
vetenskapsmännen kommer att vara fast anställda , men det kommer också att bli nödvändigt att arbeta med vetenskapsmän på konsultbasis och under dessa omständigheter är det förmodligen bättre att de , eftersom de måste resa , förflyttar sig till en central plats , där återigen parlamentets strukturer och kommissionen och rådet är baserade .
detta är min bedömning för tillfället .
det kan bli ämnet för diskussion här och annorstädes och jag kommer att lyssna på alla förslag som framläggs , men min preliminära slutsats är att denna myndighet hellre bör vara centralt placerad än i periferin .
jag befinner mig i en mycket svår position för jag kan inte ändra föredragningslistan .
jag skulle vilja föreslå att ni tar upp detta med era politiska grupper och på talmanskonferensen .
om ni känner att dessa sessioner efter ett uttalande från kommissionen är viktiga skulle jag föreslå att vi kräver mer tid än den halvtimme som är avsatt för dem .
vid detta tillfälle har vi haft sex minuter frågor från ledamöterna och 29 minuter svar från kommissionären , samt hans uttalande .
som ni ser är en halvtimme egentligen inte i närheten av vad som vore tillräckligt för en sådan sittning .
jag hoppas att ni diskuterar detta i era politiska grupper så att vi kan få en mer välstrukturerad sittning med kommissionen vid framtida tillfällen .
frågestund ( kommissionen )
nästa punkt på föredragningslistan är frågor till kommissionen ( b5-0003 / 2000 ) .
jag vill meddela att frågestunden kommer att pågå i cirka en timme och femton minuter .
vi kommer dock att begränsa tiden något , eftersom tolkarna arbetar oavbrutet under dagens sammanträde .
jag överlämnar ordet till purvis för en ordningsfråga .
jag protesterar mot att vi drar ned på tiden för frågestunden . det är ett av de få tillfällen då vanliga ledamöter har en chans att få tala och jag ber er att utöka den till en och en halv timme som på föredragningslistan .
så säger föredragningslistan och jag anser att vi skall hålla oss till den .
faktum är , käre kollega , att vi enligt föredragningslistan borde börja kl. 17.30 , och ni har klockan framför er .
jag hoppas åtminstone att sammanträdet inte fortsätter långt in på natten .
fråga nr 28 från ( h-0781 / 99 ) :
angående : anläggning av kärnkraftverk i det jordbävningsdrabbade turkiet de två senaste jordbävningarna i turkiet som båda mätte över 7 grader på richterskalan föder stor undran över att turkarna envist framhärdar med att uppföra dyra kärnkraftsreaktorer i akköy - samtidigt som energiförråden från ataturk-dammarna exporteras till tredje länder och eu gör nedskärningar i sin budget för att kunna bevilja pengar för restaureringsarbetena med anledning av de skador som jordbävningarna förorsakat .
de turkiska planerna för utvecklande av kärnkraft , som inte verkar ta hänsyn vare sig till de faror som dessa innebär för invånare eller ekosystem i turkiet och angränsande områden , föder misstankar om att det kanske bakom dessa planer döljer sig medvetna beslut , som fattats av de turkiska politiska och militära makthavarna , om att tillägna sig kärnteknik som i framtiden skall möjliggöra framställning av kärnvapen . fog för dessa misstankar finner man bland annat i det faktum att landet har för avsikt att skaffa sig reaktorer av kanadensisk typ , det vill säga likadana som de reaktorer som finns i indien och pakistan .
vilka åtgärder tänker kommissionen vidta för att kärnkraftsolyckor skall kunna undvikas och spridande av kärnvapen skall kunna hindras i ett land som önskar ansluta sig till eu och som spenderar enorma summor på program för utvecklande av kärnteknik samtidigt som det slukar europeiska medel beviljade av eu , medel som det erhåller i form av ekonomiskt bistånd ?
jag överlämnar ordet till verheugen som företrädare för kommissionen .
. ( en ) kommissionen följer med intresse det planerade bygget av ett kärnkraftsverk i akkuyu i turkiet och inser vikten av att säkerställa att det nya verkets konstruktion följer högsta internationellt godkända standard för kärnenergisäkerhet .
enligt vad vi har erfarit har inte beslutet om val av entreprenör tagits ännu .
kommissionen noterar det faktum att turkiet har undertecknat och ratificerat konventionen om kärnenergisäkerhet och att ansvaret för att bevilja tillstånd och reglera förläggning , konstruktion , igångkörning , drift och nedstängning av kärnkraftverk i turkiet helt åvilar den turkiska atomenergimyndigheten .
kommissionen har inget mandat att sätta upp gränser för beslut som fattas av något land om energiproduktion , kärnkraften inbegripen .
som kommissionär wallström berättade under utfrågningen i europaparlamentet i september 1999 kommer kommissionen att ta upp frågan om kärnenergisäkerhet och strålskydd vid alla relevanta möten med den turkiska regeringen i framtiden och det gläder mig att kunna informera er om att jag kommer att ha ett möte med den turkiske utrikesministern om några dagar och förstås kommer att ta upp frågan .
kommissionen är särkilt medveten om allmänhetens oro för den uppmätta seismiska aktiviteten i området kring ecemis-förkastningslinjen i närheten av den plats där verket föreslås bli placerat .
enligt information från internationella atomenergiorganet tar man i verkets utformning hänsyn till möjligheten av jordbävningar som är kraftigare än några som någonsin har registrerats i området och mer än tio gånger kraftigare än den som uppmättes i adana i juni 1998 .
stora utformningsmässiga marginaler skapas för att säkerställa att verket kan drivas säkert i enlighet med miljöförhållandena på platsen .
kommissionen är också medveten om oron för den möjliga avsikten att använda verket för att producera material till vapen .
den noterar det faktum att turkiet har undertecknat och ratificerat fördraget om icke spridning av kärnvapen och därefter har slutit ett omfattande avtal om garantier med internationella atomenergiorganet .
jag tackar för svaret .
jag vill göra följande påpekande : turkiet är nu kandidatland .
genom detta projekt vill landet öka sin energikapacitet med 2 procent .
samtidigt vill det förvärva reaktorer av typ cadou från canada , reaktorer som redan har använts för att framställa pakistans och indiens kärnvapen , som det har framkommit .
mot denna bakgrund finns det en mycket allvarlig risk att någon vettvilling kommer fram till att den geostrategiska balansen i kaukasus kräver att det i närheten finns ett land med kärnvapenteknik detta är den politiska aspekten .
jag övergår nu till den tekniska aspekten .
säkerhetskoefficienten vid anläggningar av detta slag - och jag talar nu som ingenjör - har inget samband med att risken för reaktorhaveri ökar 10 eller 20 gånger .
när det råder tveksamhet , använder man i dessa fall simulatorer .
vi kan emellertid inte använda simulatorer , när det gäller kärnkraft .
därför måste alla områden med hög seismisk risk a priori vara uteslutna , när det gäller kärnkraftsanläggningar av denna typ .
eftersom europeiska unionen och kommissionen nu har andra möjligheter i fråga om turkiet , bör man också diskutera vissa frågor som gäller säkerheten i området som helhet , men också frågan om turkiets fredliga utveckling i europeiska unionens sammanhang .
. ( en ) för några veckor sedan hade vi en debatt i parlamentet om kärnenergiäkerhet med speciell inriktning på kandidatländerna .
jag har förklarat kommissionens inställning .
man måste acceptera det faktum att det inte finns något regelverk i gemenskapen för kärnenergisäkerhet .
så det vi gjorde var att använda politiska medel för att övertyga vissa kandidatländer om att vi måste ha nedstängningsplaner för somliga reaktorer som inte anses möjliga att uppgradera .
i fråga om turkiet är det annorlunda .
kärnkraftverket finns inte än .
jag har redan sagt att turkiet har undertecknat icke-spridningsavtalet och konventionen om kärnenergisäkerhet .
om vi under fullbordandet av detta kärnkraftverk finner att det finns säkerhetsproblem kommer vi att diskutera detta med turkiet .
om slutsatsen är att turkiet planerar att bygga ett kärnkraftverk som inte uppfyller normala europeiska säkerthetsnormer kommer vi att göra samma sak som med litauen , slovakien och bulgarien .
herr talman ! kommissionären sade att turkiet har undertecknat icke-spridningsavtalet och kärnenergisäkerhetsfördragen : varför skulle det finnas något som helst tvivel på att turkiets kärnkraftverk inte skulle bli precis lika säkert som något annat i gemenskapen , och skulle kommissionären vara beredd att inta en något mer kraftfull ståndpunkt mot souladakis i denna fråga ?
. ( en ) jag anser att en parlamentsledamot har rätt att ta upp det han oroar sig och är rädd för .
jag är inte orolig för detta .
jag tror att turkiet till fullo godtar normerna och kriterierna i konventionen om kärnenergisäkerhet och i icke-spridningsavtalet , men det finns otvivelaktigt en oro bland allmänheten i europa och jag tycker att det är helt rätt att diskutera den här i parlamentet .
fråga nr 29 från ( h-0786 / 99 ) :
angående : vapen med utarmat uran har kommissionen gjort några utredningar av hur staterna inom eu kan komma att påverkas av gränsöverskridande föroreningar som uppstått till följd av att det i kosovokonflikten använts vapen med utarmat uran ?
om inte : varför inte ?
härmed överlämnar jag ordet till wallström , som företrädare för kommissionen .
. ( en ) tack för er fråga , herr bowe .
europeiska kommissionen har övervakat konfliktens miljökonsekvenser från det att natoaktionen inleddes .
redan i juni förra året finansierade kommissionen en första utredning .
den genomfördes av det regionala utvecklingscentrumet för central- och östeuropa och slutsatsen var att ingen storskalig ekologisk katastrof hade ägt rum .
denna första bedömning har inte ändrats av senare bevis eller analyser .
kommissionen har också varit intimt inblandad i framtagandet av den rapport som nyligen utgavs av förenta nationernas miljöprogram - insatsstyrkan på balkan .
detta är den hittills mest detaljerade och omfattande rapporten om kosovokrigets miljökonsekvenser och jag rekommenderar dem av er som ännu inte har tagit del av den att göra det .
användningen av utarmade uranvapen var en av de många frågor som behandlades och denna rapport finns nu lätt tillgänglig , också på internet .
insatsstyrkan på balkan hindrades av det faktum att det praktiskt taget inte fanns någon information om den faktiska användningen av dessa vapen under kriget .
på sin faktainsamlingsresa fann de inga tecken på kontamination i kosovo .
detta utesluter dock inte att områden i kosovo kan vara kontaminerade med utarmat uranium .
av en skrivbordsutvärdering tillsammans med en faktainsamlingsresa dras i rapporten slutsatsen att eventuella risker begränsas till ett område kring målet .
framtida åtgärder kommer att genomföras inom ramen för stabilitetspakten för sydöstra europa .
en särskild regional plan för rekonstruktion av miljön håller också på att tas fram .
den kommer att bilda ramen för nödinsatser för att bekämpa krigsskador , om sådana skulle behövas .
herr talman ! först av allt ber jag att få tacka kommissionären för detta mycket matnyttiga svar .
det är tydligt att kommissionen har övervägt detta problem , och jag är glad att man i de rapporter som hittills har framtagits granskar frågan ingående .
men jag skulle vilja påpeka att oron för utarmade uranvapen gäller sättet de används på .
detta uranium blir luftburet och man andas in det . det skulle nu faktiskt kunna vara så att delar av befolkningen i kosovo bär på detta , med mycket mer långsiktiga effekter än man hittills kunnat fastställa .
detta verkar vara det händelsemönster som har framkommit efter användningen av utarmade uranvapen i gulfkriget .
jag skulle därför vilja fråga kommissionen om den skulle vilja överväga att fortsätta övervakningen och under hur lång tid de skulle kunna tänka sig att i framtiden övervaka för att se vilka de långsiktiga konsekvenserna blir , inte bara av utarmade uranvapen utan också en del av de andra miljökonsekvenser vi vet har uppstått åtminstone lokalt i kosovo ?
hur länge kommer ni att fortsätta att utvärdera konsekvenserna av dessa vapen ?
. ( en ) tack för den frågan , herr bowe .
vi måste återigen hävda att det fortfarande inte är bekräftat att utarmat uran användes i kriget och att inget utarmat uran har upptäckts under upprensningen i kosovo .
men de symptom och de problem ni nämnde kan finnas där , och de kan vara konsekvenser av användningen av utarmat uran .
detta nämns också i rapporten .
inga gränsöverskridande konsekvenser har upptäckts och de flesta vapnen måste ha använts inom förbundsrepubliken jugoslaviens territorium .
problemet är att landets nuvarande politiska isolering innebär att tillträdet till detta område är begränsat .
förenta nationerna har ett stort ansvar , för denna rapport vänder sig till dem , så de måste ta sitt ansvar .
men genom denna regionala och miljömässiga rekonstruktionsplan kan vi fortsätta övervakningen och det bistånd vi kan ge och detta är , för närvarande , den slags ram vi kan använda för europeiska unionens arbete .
uppföljning är viktig och den ger medlemsstaterna , liksom förenta nationerna och kommissionen , någonting att tänka på när den handlar om militära hemligheter och deras konsekvenser för miljön .
den har också en långsiktig påverkan på tänkandet när det gäller användningen av detta slags vapen .
herr talman , fru kommissionär ! om några månader kommer återigen hundratusentals semesterfirare att fara till den adriatiska kusten och tillbringa sin sommarledighet där .
som vi känner till från nyhetsrapporterna , har bomber och vapen fällts i närheten av kusten .
kan ni bekräfta att semesterfirarna denna sommar kan bada riskfritt i adriatiska havet , och har man planerat åtgärder för att undersöka hur hotbilden ser ut ?
. ( en ) jag önskar att jag kunde garantera mycket , men tyvärr kan jag inte det .
vi gör våra bedömningar utifrån rapporter som denna och de sändebud vi skickar ut för att kontrollera sådana här saker .
det är detta vi grundar oss på när vi råder människor vad de skall göra .
det vi har sett är att krig påverkar miljön på lång sikt och detta är farligt .
på miljöområdet har vi just antagit ett direktiv om föroreningar till havs .
detta innefattar kulor och vapen och så vidare och är ett förvarningssystem .
tyvärr kan vi inte utfärda garantier utan bara fortsätta att övervaka och försöka genomföra upprensningar .
jag ville fråga kommissionären om det är sant att soldater från natos väpnade styrkor som nu är stationerade i denna region genomgår särskilda kärnstrålningskontroller och att samma åtgärder inte tillämpas på civilbefolkningen i området ?
. ( en ) jag kan inte svara på den frågan .
jag har inte all den information som fordras för att svara ordentligt när det handlar om läkarkontroller och så vidare .
vad vi vet från miljösidan är det jag redan har nämnt , att det nu finns en plan för rekonstruktion av miljön , men när det gäller läkarkontroller har jag ingen information .
jag kan naturligtvis gå tillbaka och se om vi kan hitta den information som behövs .
fråga nr 30 från ( h-0793 / 99 ) :
angående : utnämning av ett särskilt eu-sändebud för tibet för 1998 registrerade den tibetanska exilregeringen att över 4 000 tibetaner flytt över himalayabergen till friheten med fara för liv och lem .
många av flyktingarna drabbades därvid av allvarliga förfrysningsskador och många dog .
den tvärpolitiska gruppen &quot; tibet &quot; är mycket bekymrad över den allt värre situationen i tibet och det står klart att europeiska unionens nuvarande politik inte räcker till för att uppnå resultat vad gäller de svåra kränkningar av de mänskliga rättigheterna som tibetanerna i tibet utsätts för varje dag .
den tvärpolitiska gruppen &quot; tibet &quot; , som verkligen oroar sig över de fortsatta kränkningarna av de mänskliga rättigheterna i tibet och önskar stödja dalai lamas förslag om en dialog med den kinesiska regeringen för att lösa situationen i tibet , uppmanar därför kommissionen att utnämna ett särskilt sändebud för tibet , som skall sköta europeiska unionens angelägenheter i denna fråga och bemöda sig om att föra samman tibetanska och kinesiska företrädare och / eller myndigheter i en dialog .
när kommer kommissionen att utnämna ett särskilt sändebud för tibet ?
jag överlämnar ordet till patten , som företrädare för kommissionen .
. ( en ) den oro europaparlamentet uttrycker för tibet delas av många .
jag har länge trott på behovet att bestämt och rättframt för de kinesiska myndigheterna framhålla vår inställning i frågor om mänskliga rättigheter också i tibet .
europeiska unionen gjorde detta vid toppmötet mellan europeiska unionen och kina förra månaden och pressade kineserna i ett antal frågor om mänskliga rättigheter , däribland tibet .
vi uppmanade åter kina att inleda en dialog med dalai lama .
jag uppmanar igen kina att göra det .
vi kommer att fortsätta att ta upp tibet med de kinesiska myndigheterna .
vi gör också en del andra saker : inom dialogen mellan europeiska unionen och kina om mänskliga rättigheter har vi inriktat oss på ett antal praktiska steg , däribland att skicka ut experter på uppdrag till tibet , planera program för utvecklingsbistånd och verksamhet inom hälsa och utbildning för tibetanerna .
utnämningen av ett särskilt eu-sändebud för tibet skulle främst vara en fråga för rådet att besluta om och parlamentet kanske vill ta upp frågan direkt med dem .
men för egen del är jag inte säker på att det skulle bidra så mycket till våra ansträngningar i praktiken .
det skulle troligen inte ha någon större inverkan på de kinesiska myndigheterna och vi har redan effektiva kommunikationskanaler med exiltibetanerna .
jag tycker också att det är angeläget att akta sig för en exponentiell ökning av särskilda sändebud , hur gott syftet än är .
herr talman , herr patten ! ni har naturligtvis utmärkta erfarenheter på grund av ni levt i kina , och ni vet mycket väl hur tibetanerna anstränger sig för att åstadkomma en dialog , vilket hittills alltid har förhindrats .
men om ert svar blir att vi skall vända oss till &quot; mister gusp &quot; , alltså till solana , då befarar jag att det är en ensidig inriktning av utrikespolitiken .
er ansats , som jag mycket väl rekommenderar som en sammanhållande ansats , har ju inspirerats av de mänskliga rättigheterna ; jag håller helt med om att vi måste ta oss an frågan om human rights .
anhållandena , tortyren , stympningen av unga kvinnor och liknande , det är ju absolut diskussionsämnen som man kan ägna sig åt en hel kväll .
om vi inskränker det och säger att rådet här också är ansvarigt , så befarar jag att dessa frågor om de mänskliga rättigheterna inte kommer i dagen tydligt nog .
möjligheten att å ena sidan betona ekonomi och handel , men att mycket väl integrera de mänskliga rättigheterna , vore en åtgärd där vi egentligen satsar på kommissionens partnerskap , och inte säger att det är en fråga för rådet .
. ( en ) låt mig klargöra för er vilken inställningen är .
jag sade ingenting annat än sanningen när jag sade att utnämningen av särskilda sändebud är en fråga för rådet .
det råkar vara så att vi hanterar de budgetmässiga konsekvenserna och rådet utser vederbörande .
somliga kanske tycker att denna budgetfråga borde ses över på sikt .
om vi lämnar det , för sådant är läget , innebär inte detta att vi inte har en åsikt och en befogenhet i fråga om mänskliga rättigheter , jag hoppas väldigt mycket att kommissionen under de närmaste månaderna kommer att kunna ta fram ett meddelande om mänskliga rättigheter där vi bland annat påpekar att det inte finns någon som helst motsättning mellan en omsorg om mänskliga rättigheter i kina eller på andra håll i världen och europeiska unionens handelsmässiga , kommersiella och andra intressen .
jag har länge ansett att vi alla bör erkänna att de länder som det är bäst att göra affärer med är de länder som behandlar sina egna medborgare mest anständigt - överallt i världen .
jag upprepar att vi har framfört vår uppfattning om tibet till kina .
under de få månader som jag har varit kommissionär har det hänt två gånger , först i new york vid vårt möte med minister tang och nyligen vid mötet i peking och vi kommer att fortsätta att ge uttryck för denna oro .
om jag får rekommendera en bok till er , eftersom jag inser att ni är intresserad av dessa frågor , rekommenderar jag en bok om tibet som gavs ut precis innan jul och som är skriven av den framstående journalisten isabel hilton .
herr talman ! jag vill börja min tilläggsfråga med den tibetanska hälsningen , som betyder lycka och fred .
i tibet handlar det inte bara om de mänskliga rättigheterna och miljön , utan det handlar om ett unikt kulturarv , som också kan förmedla viktiga värden till oss européer , exempelvis ro , stillhet , medkänsla , compassion , som dalai lama säger .
frågan är nu vad kommissionen kan göra för att på ett mer konkret sätt stödja hans helighet dalai lama och hans förslag till en fredlig lösning av tibet-frågan ?
jag vill påpeka att om man inte gör någonting kommer det att leda till att den tibetanska kulturen dör ut och att det tibetanska folket försvinner .
. ( en ) jag känner stor sympati för vad ni sade om kulturarv och om den buddhistiska traditionen .
liksom ni har jag läst dalai lamas självbiografi .
det är en mycket rörande berättelse , inte bara om hans skyldigheter i och gentemot tibet utan också om hans andliga åskådning .
kommissionen har , liksom andra , uppmanat till dialog .
dalai lama har gjort klart att han önskar en fredlig dialog .
jag önskar att de kinesiska myndigheterna hade svarat konsekvent och positivt på denna invit från dalai lama .
vid eller omkring tiden för president clintons besök i kina gav presidenten i folkrepubliken kina intryck av att dialog stod på dagordningen .
det skulle vara mycket välgörande , inte bara för tibet och för alla de som tror på fred och stabilitet i asien , utan det skulle också verkligen vara till heder för folkrepubliken kinas regering om den skulle svara på dessa försök att inleda en dialog .
fråga nr 31 från ( h-0795 / 99 ) :
angående : stadgan om god förvaltning inom eu som avvisats av kommissionen enligt uppgifter i pressen har kommissionen avvisat det förslag om medborgarnas rätt till god förvaltning inom eu , vilket framlagts av den europeiska ombudsmannen jacob söderman .
kommissionen har själv godkänt tanken på en stadga för god förvaltning men kom nu att avvisa det detaljerade förslaget och framlade i stället en rad kompletterande föreskrifter om bättre service .
stämmer de ovannämnda uppgifterna ?
vad finns det för orsak till att kommissionen handlat som den gjort och hur vill kommissionen förklara den skillnad mellan ord och handling som på det här viset uppstått på tal om förnyandet av eu : s förvaltning ?
tycker kommissionen att det inträffade stämmer överens med det fempunktsprogram som europaparlamentet och kommissionen kom överens om i september och är kommissionen beredd att framlägga ett detaljerat förslag till en stadga för god förvaltning i sådan form att också parlamentet har en möjlighet att ta ställning till det ?
. ( en ) den tidningsartikel som ni hänvisar till tycks mig vilseledande och felaktig .
i november 1999 antog kommissionen vid förstabehandling en uppförandekod för tjänstemännen som skulle införlivas med arbetsordningen .
för närvarande rådgör kommissionen med sina tjänstemannarepresentanter om detta dokument , och denna process kommer att slutföras under de närmaste veckorna .
kommissionen kommer då att anta koden vid andrabehandling .
man bör notera att den nya kommissionen på eget initiativ omedelbart följde upp den europeiske ombudsmannens beslut från 28 juli 1999 i hans utredning om koden .
kommissionen skulle speciellt vilja betona att vi när vi upprättade denna kod har anammat alla ombudsmannens förslag till rekommendationer .
koden kommer att bli ett dokument som uteslutande handlar om kommissionens tjänstemäns förhållande till allmänheten .
den kommer att antas genom ett juridiskt bindande beslut i kommissionen som kommer att offentliggöras i europeiska gemenskapernas officiella tidning .
dokumentet har sammanställts med full hänsyn till de bestämmelser som finns i det förslag som den europeiske ombudsmannens kontor har upprättat .
enligt bestämmelser i fördragen om detta är det kommissionen själv som ansvarar för att fastställa sin arbetsordning .
det är emellertid självklart att kommissionen håller fast vid principen om regelbunden politisk dialog med europaparlamentet om alla aspekter av administrativa reformer .
herr talman ! jag vill tacka kommissionären .
jag frågar ändå , när är det meningen att denna stadga äntligen skall träda i kraft ? med tanke på att den har hållit på att utarbetas ända sedan 1997 .
. ( en ) tidningsartiklarna var vilseledande .
jag tror inte att det finns någon skillnad mellan oss och ombudsmannen .
det finns en fråga om den rättsliga grunden och där har vi inhämtat råd och jag tror att vi har väl på fötterna där .
jag vill upprepa att ledamöter som liksom den ledamot som ställde frågan är speciellt intresserade av denna fråga säkert vill föra en dialog om den .
det är ytterst viktigt och jag förstår er oro .
jag vill tacka kommissionen för det som jag uppfattar som ett mycket positivt svar .
för säkerhets skull skulle jag vilja ha en bekräftelse på att det verkligen är så , att det inte finns någon del av jacob södermans förslag , vad gäller kommissionen och den goda förvaltningen , som kommissionen tycker är oacceptabel .
är det korrekt att alla delar av förslaget kommer att godtas till sitt innehåll ?
. ( en ) låt mig läsa vad det står i mitt sammandrag - och eftersom det står där måste det vara sant !
&quot; jag skulle återigen vilja betona att kommissionen har godtagit alla ombudsmannens rekommendationer i hans förslag till rekommendationer från juli 1999 &quot; .
båda dokumenten , det vill säga kommissionens dokument och ombudsmannens förslag , täcker i stort sett samma saker .
den enda substantiella fråga som har uppstått är den rättsliga grunden .
jag kan gå in på den i detalj om ni vill men det finns inget tvivel om att vi är ense med ombudsmannen i denna viktiga fråga .
vi tar gärna med pattens kommentarer i vår litteraturförteckning , som ett komplement till ledamöternas favoritlektyr .
eftersom frågeställaren är frånvarande , bortfaller fråga nr 32 .
jag ber vitorino om ursäkt för parlamentets ohövliga agerande , vilket jag beklagar .
enligt arbetsordningen har parlamentet ingen skyldighet att svara .
jag önskar er en fortsatt bra dag .
frågor till nielson som har ersatts av patten
frågorna 33 och 34 i andra delen av frågor till kommissionen är riktade till nielson .
nielson kan inte närvara här i dag , eftersom han befinner sig i sydafrika .
jag kan meddela att kommissionens vice ordförande loyola de palacio har skickat ett brev där hon förklarar detta och meddelar att patten kommer att vara den som besvarar dessa frågor .
fråga nr 33 från ( h-0829 / 99 ) :
angående : mainstreaming i eu-biståndet ministerrådet utarbetade redan 1995 riktlinjer för integrering av ett jämställdhetstänkande ( mainstreaming ) i hela eu : s biståndspolitik .
riktlinjerna kräver att all personal som arbetar med utvecklingsfrågor skall få kontinuerlig fortbildning i &quot; gender mainstreaming &quot; , men under de senaste åren har bara ett 50-tal personer utbildats och fortfarande finns ingen obligatorisk jämställdhetsutbildning på generaldirektoratet för bistånd .
att låta ett jämställdhetstänkande genomsyra den totala verksamheten ( mainstreaming ) innebär att hänsynen till jämställdhet mellan kvinnor och män ingår som en självklar del i alla former av utvecklingspolicy , strategier och insatser .
för att möjliggöra detta måste rådets riktlinjer om mainstreaming tillämpas i sin helhet .
nuvarande personal måste få obligatorisk utbildning i jämställdhetsfrågor och 1-2 dagars utbildning i jämställdhetsfrågor bör ingå som en nödvändig del i generaldirektoratet för bistånds obligatoriska introduktionskurser för nyanställda .
är kommissionen beredd att vidta dessa åtgärder ?
. ( en ) får jag först av allt betona hur ledsen min kollega nielson var att han inte kunde vara här , men ni som bryr er om dessa utvecklingsfrågor vet säkert hur viktigt hans uppdrag är , att försöka se till att vårt avtal med sydafrika överlever .
kommissionen är beredd att titta på möjligheterna att göra en genomgång av jämställdhets- och utvecklingsfrågor till en del av de så kallade introduktionskurserna för ny personal , någonting som redan har förekommit , fast inte regelbundet får jag erkänna .
utbildning av personal som flyttar till delegationerna i de olika regionerna är en annan inkörsport .
utbildningen skulle då genomföras automatiskt utan att vara obligatorisk .
vi siktar också på att lägga in utbildning i dessa frågor i den grundkurs i projektadministration våra tjänstemän genomgår .
vi vill att detta slags utbildning så långt som möjligt skall vara automatiskt inbyggd i programmen från början i stället för att man skall hantera den separat senare .
min personliga inställning som före detta utvecklingsminister är att dessa frågor själva borde integreras och tacklas som en del av utbildningen , inte göras till något slags frivilligt tillval .
strävan efter jämställdhet skall på alla nivåer genomsyra arbetet vid generaldirektoratet för bistånd .
den skall inte tillföras som &quot; något vid sidan om &quot; .
detta måste naturligtvis leda till en omformulering av utvecklingsmål och strategier samt en omvandling av institutioner och processer , så att såväl kvinnors som mäns prioriteringar och behov avspeglas på ett bättre sätt .
vidare måste åtgärder mot könsgrundade skillnader vidtas .
jämställdhet måste genomsyra inte bara projekt och program , utan också alla övergripande mål , handlingsplaner och strategier .
det ser ut som om vi är överens om detta .
men ansvaret för att vederbörlig uppmärksamhet ägnas jämställdhet ligger hos avdelnings- och enhetschefer .
om inte cheferna besitter den professionella kompetens som krävs , så sker ingenting - gender mainstreaming bortprioriteras .
ytterst få i ledningen av generaldirektoratet för bistånd , dvs. enhetschefer och ännu högre chefer , har deltagit i de genderkurser som har anordnats .
endast en chef har deltagit i genderutbildningen en halv dag .
vad är kommissionen beredd att göra för att se till att enhetschefer och chefer på ännu högre nivå genomgår nödvändig genderutbildning ?
det har hänt att gender har ingått i den obligatoriska introduktionskursen för nyanställda , men då bara en till två timmar per kurs .
detta begränsade utbildningsmoment har dock strukits från alla introduktionskurser som har ägt rum under senare tid .
som jag i min fråga påpekar , krävs det inte att en till två timmar , utan att en till två dagar ägnas åt ämnet .
min fråga är : är kommissionen verkligen beredd att fullfölja de antagna riktlinjerna för gender mainstreaming på generaldirektoratet för bistånd ?
. ( en ) jag tar verkligen frågan om integrering av ett jämställdhetsperspektiv på allvar , och det gör min kollega kommissionär nielson också .
jag skall inte tjata om böcker , men jag har just läst en bok av david landis barnhill om vad det är som gör att vissa länder blomstrar och andra inte , och det är intressant att se den betydelse han fäster vid jämställdhetsfrågor för ekonomisk framgång och politisk stabilitet i olika samhällen under årtusendena .
för det andra anser jag att även om den utbildning vi talar om inte bör vara obligatorisk - när allt kommer omkring finns ingen obligatorisk utbildning om någonting hos kommissionen - bör den vara väsentlig .
och eftersom den bör vara väsentlig skulle man hoppas att alla skulle se till att de hade tillräcklig jämställdhetsutbildning .
det gäller alla , på alla nivåer .
det är inte någonting som högre tjänstemän skall bedöma som lämpligt för sina underställda , men tro att de själva är för vuxna eller för högt uppsatta för att genomgå .
för det tredje är ett av de bästa sätten att angripa denna fråga att integrera jämställdheten som en viktig och gränsöverskridande fråga i de mest populära kurserna för utvecklingstjänstemän och framför allt kanske i kursen om projektadministration som är nyckeln till god administration av projekt på fältet .
så jag håller till stor del med om det ni sade .
jag hoppas att det angreppssätt vi har anammat visar på både ett praktiskt sinnelag och vikten av att detta får den uppmärksamhet det förtjänar .
. ( en ) sedan 1991 ger gemenskapen ett betydande ekonomiskt stöd till de nya oberoende staterna och däribland länderna i centralasien .
större delen av europeiska unionens stöd har tillhandahållits inom ramen för tacis-programmet .
1998 och 1999 erhöll kirgizistan , kazakstan , uzbekistan och turkmenistan tekniskt bistånd på 75 miljoner euro .
detta bistånd har gagnat alla områden , särskilt jordbruket , infrastrukturutvecklingen , privatekonomin och stärkandet av institutionerna .
tadzjikistan har av säkerhetsskäl inte kunnat dra nytta av tacis fullt ut , men ett återuppbyggnadsprogram på 7,2 miljoner euro har funnits på plats under 1998 och 1999 .
förutom de nationella programmen har europeiska unionen stött viktig regional verksamhet inom energi- , transport- och miljösektorerna .
livsmedelssäkerhetsprogram i centralasien inleddes 1996 efter att europeiska unionen under två år levererat livsmedelsstöd in natura .
dessa program har gagnat kirgizistan och i mer begränsad omfattning tadzjikistan .
avsatta medel för de icke-statliga organisationernas program i tadzjikistan uppgick till 7,42 miljoner euro 1998 och 1999 .
under samma period fick kirgizistan 17 miljoner euro .
sedan 1993 har kommissionens europeiska gemenskapernas kontor för humanitärt bistånd , echo , aktivt stött de mest utsatta grupperna och sektorerna i tadzjikistan och kirgizistan .
för 1998 och 1999 avsattes 3,8 miljoner euro till kirgizistan och tadzjikistan erhöll över 35 miljoner euro , huvudsakligen för livsmedel , läkemedel , vatten och hygien .
det har framgått av regelbundet återkommande utvärderingar och lägesbedömningar att europeiska unionens stöd bidrar till dessa länders stabilitet och därmed till den pågående fredsprocessen .
herr talman , herr kommissionär ! centralasien och kaspiska havet hotar ju att bli 2000-talets balkan .
därför hänger det mycket på en stabilisering av just de stora staterna turkmenistan och uzbekistan .
jag vill därför fråga er , och detta ligger ju inom ert eget ansvarsområde , hur förhandlingarna beträffande partnerskapsavtalet med dessa båda länder går , alltså de politiska förbindelserna .
det är ju direkt ert område ; min andra fråga gäller kollegan nielsens område : hur går det ekologiska samarbetet , i synnerhet beträffande vattnet och problematiken med monokulturerna av bomull , som leder till stor uttorkning .
. ( en ) under toppmötet i istanbul för några veckor sedan hade vi tillfälle att träffa och föra diskussioner med några av de centralasiatiska republikerna .
jag är mycket mån om att vi stärker våra relationer med dem .
om ni vill kan jag skicka er en detaljerad sammanställning av exakt var vi befinner oss i förhandlingarna om partnerskap och samarbetsavtal med var och en av de centralasiatiska republikerna .
alla hoppas naturligtvis att denna förutsägelse om vad som kan hända i framtiden är för pessimistisk .
men jag tvivlar inte alls på att ni har rätt när ni betonar centralasiens strategiska betydelse .
jag har tidigare hört er tala om kaukasus också .
ni har helt rätt i att en union som talar om att förhindra konflikter borde titta på vad den kan göra i dessa speciella områden för att tillse att den typ av konflikt inte uppstår som den på balkan som har orsakat så mycket förödelse och som har kostat oss en hel del mer än vi kanske skulle ha gjort av med annars , om vi hade vidtagit fler förebyggande åtgärder , om dessa hade varit möjliga .
så era kommentarer om dessa regioners strategiska betydelse är ytterst välfunna .
vi bidrar till program i regionen som har viss miljöpåverkan .
våra livsmedelsprogram hänger direkt samman med strukturella jordbruksreformer liksom med lindrande av fattigdom .
dessa program syftar i sig till att säkerställa att jordbruket får en sundare bas i dessa samhällen och inte bara går ut på att våldta jorden .
det finns en ekologisk aspekt som vi bör fortsätta att prioritera .
lägg märke till att den ledamot som ställde frågan applåderade kommissionärens svar .
det sker inte så ofta .
och dessutom har kommissionären i det här fallet inte nämnt litteraturförteckningen .
tack så mycket , herr patten , för era inlägg i dag .
fråga nr 35 från ( h-0778 / 99 ) :
angående : greklands åtgärdsplan för sysselsättningen enligt vad som framkommit vid utvärderingen av åtgärdsplanerna för sysselsättning har kommissionens kritik huvudsakligen riktats mot grekland och italien för att dessa inte på vederbörligt sätt genomfört sysselsättningspolitiken och stödåtgärderna för sysselsättningen .
i rapporten konstateras det att varken grekland eller italien ännu nått målen för förbättrad anställbarhet och att det är tvivel underkastat om den politik som avses genomföras kommer att göra det möjligt att följa riktlinjerna för hur långtidsarbetslösheten skall förebyggas eller hanteras .
i rapporten ingår också en kommentar om att grekland inte planerat några åtgärder på medellång eller lång sikt för att sänka arbetsgivarens skatter och försäkringsavgifter i samband med anställande och att det dessutom inte föreligger några exakta siffror över sysselsättningen .
kan kommissionen upplysa om greklands regering ingått några särskilda åtaganden för hur problemet med ungdoms- och långtidsarbetslöshet kunde angripas och vilka dessa åtaganden i så fall är ?
har regeringen lagstiftat om och infört något system för hur växlingarna i sysselsättning skall kunna fastställas , registreras och övervakas eller handlar merparten åtgärder fortfarande bara om att räkna dem som är utan arbete ?
som svar på papayannakis fråga kan jag säga att det i åtgärdspaketet för sysselsättning 1999 framförde kommissionen vissa förslag och rekommendationer till grekland i syfte att effektivisera sysselsättningsåtgärderna .
den viktigaste punkten var att man måste anstränga sig för att reformera den offentliga förvaltningen , där det finns problem . man måste förbättra systemet för statistisk uppföljning och vidta förebyggande politiska åtgärder i enlighet med riktlinjerna 1 och 2 i sysselsättningspaketet .
jag måste tala om att den grekiska regeringen , inom ramen för sin arbetslöshetspolitik , har två konkreta program för 1999 : &quot; ja till yrkeslivet &quot; och &quot; tillbaka till arbetet &quot; .
jag har ännu inte fått veta det slutliga resultatet av dessa program , så att jag kan se om de kvantitativa målen har uppnåtts .
den grekiska regeringen är i dag medveten om problemet med att man inte kan registrera flödet av arbetskraft till och från sysselsättning och har därför åtagit sig , för det första , att omorganisera landets arbetsmarknadsmyndigheter , för det andra , att skapa effektiva centra för främjande av sysselsättning - detta program har redan inletts men har ännu inte avslutats - för det tredje , att införa ett lämpligt system för elektronisk registrering av sysselsättningen för att kunna följa upp alla dessa praktiska åtgärder .
i det nya programmet för perioden 2000-2006 , som finansieras av europeiska socialfonden , bör man , även med kommissionens stöd , utnyttja alla nödvändiga resurser och politiska åtgärder för att förverkliga de mål jag tidigare nämnde .
kommissionen kommer att noga följa hur den grekiska regeringen fullföljer sina åtaganden .
jag tackar kommissionsledamoten för hennes svar . men , fru kommissionär , vi befinner oss i följande situation .
i fråga om arbetslöshetens omfattning ligger vi på andra plats i europa , dvs. 11,3 procent - vilket vi inte gjorde tidigare - , vi har den största ökningen av arbetslösheten , vi lägger ut minst pengar på de arbetslösa , dvs. mindre än 1 procent av bnp , medan andra länder spenderar 3-4 procent ( t.ex. frankrike , belgien och tyskland ) , och det är inte klart hur man har använt de pengar som europeiska socialfonden betalat ut , bl.a. för att bekämpa arbetslösheten .
ni säger att kommissionen har lämnat vissa rekommendationer .
jag gläder mig över detta och hoppas att man följer rekommendationerna .
men jag har väldigt länge burit på en fråga : hur har det gått med de tidigare politiska åtgärderna ?
är det någon som fått ett arbete ?
hur många har fått arbete ?
i fjol och i förfjol , om ni inte kan säga hur det är i år .
hur har det gått med yrkesutbildningen ?
dessa så omtalade utbildningscentra , är de till för att ge arbete åt dem som utbildar eller åt dem som utbildas ?
har vi några siffror ?
har vi således någon möjlighet att kontrollera hur den grekiska regeringen sköter denna politik ?
herr papayannakis ! vad jag skulle kunna svara är att vad den grekiska regeringen verkligen bör satsa på är den elektroniska statistiska registreringen av befintliga strukturer , så att de pågående programmen kan ge de kvantitativa resultat som ni talar om , men också för att möjliggöra en uppföljning som ger underlag för den politik som bör föras .
grekland har uppvisat en ökad sysselsättningsgrad och - efter vad jag kan se här - också en ökad produktivitet .
det kommissionen kan påverka är de konkreta riktlinjerna .
som ni vet , är det 22 riktlinjer som varje land bedöms efter .
de gäller tillgång till yrkesutbildning och de speciella åtgärderna för långtidsarbetslösa .
i fråga om alla dessa riktlinjer kommer kommissionen att försöka få fram kvantifierbara data och konkreta uppgifter om förverkligandet av gemenskapens riktlinjer för perioden 2000-2006 .
fråga nr 36 från ( h-0782 / 99 ) :
angående : det danska systemet för förtidspension har kommissionen godkänt det danska systemet för förtidspension i sin helhet ? råder det eventuell oenighet mellan danmark och kommissionen på andra socialpolitiska områden ?
det danska pensionssystemet , eftarløn , innebär att pension endast kan utgå till dem som är bosatta i danmark och till dem som uppfyller kravet på att ha arbetat en viss tid i detta land .
det finns arbetstagare som framfört klagomål till europeiska kommissionen för att de inte har rätt till pension .
de danska myndigheterna anser inte att gemenskapslagstiftningen tvingar dem att betala ut denna ersättning till förtidspensionerade arbetstagare , när dessa inte uppfyller villkoren enligt dansk lag .
det bör noteras att gällande förordning om socialförsäkringssystem för närvarande inte omfattar några bestämmelser om förtidspensionering , och kommissionen har föreslagit vissa förändringar i förordningen , vilka emellertid ännu inte har avgjorts av rådet .
eg-domstolen har hittills ännu inte tagit ställning till eftarløn , men man skulle på goda grunder kunna hävda att bosättningsvillkoren inte är förenliga med de allmänna kraven på förbud mot diskriminering på grund av medborgarskap .
europeiska kommissionens tjänsteenheter har inlett ett förfarande med möten och överläggningar med den danska regeringen för att kunna nå fram till en gemensam lösning .
det senaste mötet i denna fråga hölls i november 1999 , och vi avvaktar slutliga förslag från kommissionens tjänsteenheter om huruvida det kan bli aktuellt med ett ingripande mot danmark .
jag lade märke till att kommissionsledamoten inte gav något direkt svar på frågan om det danska förtidspensioneringssystemet i sin helhet är godkänt av kommissionen , men det framgick ju indirekt att svaret var nekande .
jag vill be kommissionsledamoten att uttryckligen bekräfta att systemet inte är godkänt av kommissionen .
kommissionen gjorde ju mer än bara antydde att man starkt överväger att ta upp hela frågan om det danska förtidspensioneringssystemet i domstolen i luxemburg , just med den utgångspunkt att det här föreligger en faktisk diskriminering i förhållande till icke-danska arbetstagare som inte kan uppfylla villkoren till följd av att de inte arbetat under den tidsperiod som krävs enligt det danska systemet .
jag vill fråga kommissionären om hon kan ange några ungefärliga tidsperioder i detta sammanhang , eftersom det är ett problem som måste få ett avgörande i den danska socialpolitiska debatten .
jag skulle alltså vara tacksam om kommissionären skulle kunna utveckla denna fråga .
herr parlamentsledamot ! vad jag skulle vilja framhålla är att det såväl i danmark som i många andra länder finns problem i fråga om tolkningen av direktiven , när de skall införlivas med respektive lands lagstiftning .
detta är ett sådant fall. och det pågår en diskussion mellan den danska regeringen och kommissionen , för att frågan skall kunna lösas på bästa sätt , till gagn för de arbetstagare som uppfyller villkoren och som , enligt gällande lagstiftning , har denna rätt till pension .
för att bara helt kort knyta an till den sista punkten . jag uppmanar kommissionen att göra det helt klart att kommissionens invändningar , för vad de är värda , inte på något sätt skulle inkräkta på danska medborgares rätt att dra nytta av denna plan utan att kommissionen bara är angelägen , vilket den har rätt att vara enligt gemenskapens lagar , om att säkerställa att planen gäller alla gemenskapsmedborgare som uppfyller villkoren .
jag anser att svaret är kort och tydligt .
det är naturligtvis så som ni sade .
det kommer inte att bli något problem med de danska medborgarna , och det är inte där problemet ligger .
problemet gäller danska eller andra medborgare , som är bosatta utanför danmark .
fråga nr 37 från ( h-0791 / 99 ) :
angående : arbetstidsdirektivet sjukhusläkare , som inte är konsulterande , omfattas inte av arbetstidsdirektivet från 1993 och inte heller av förslaget till ändring av rådets direktiv ( kom ( 98 ) 0662 - c4-0715 / 98-98 / 0318 ( syn ) ) . vilka åtgärder föreslår kommissionen för att säkerställa att skyddsnivån för dessa läkare är jämförbar med den som fastställs i direktivet från 1993 ?
fråga nr 38 från ( h-0805 / 99 ) :
angående : åtgärder för att öka jämställdheten mellan könen en av de arbetsgrupper av kommissionsledamöter som har aviserats av ordförande prodi har som mål att främja åtgärder för ökad jämställdhet mellan könen ( införlivande av jämställdhetsaspekten , så kallad mainstreaming ) .
vilka kommissionsledamöter ingår i denna grupp ?
hur många gånger har de träffats hittills ?
vilka konkreta åtgärder har diskuterats ?
frågan innehåller flera delfrågor .
den gäller kommissionens särskilda kommitté som sysslar med jämställdhetsfrågor .
de kommissionsledamöter som medverkar är ordföranden prodi , vice ordföranden kinnock , reading och jag själv .
kommitténs sammanträden är öppna , och det första sammanträdet hölls den 11 januari 2000 .
vi diskuterade tre allvarliga frågor : den första gällde det femte kvinnoprogrammet , som vi efter min föredragning hade en första diskussion om , den andra gällde busquins rapport om undersökningen av kvinnors deltagande i forskning och vetenskap , och den tredje gällde kinnock , som informerade kommissionen om ansträngningarna att ta hänsyn till jämställdhetsaspekten i det omfattande reformarbete som i dag pågår inom gemenskapen .
tack för ert svar , fru kommissionär , men jag måste beklaga att det dröjde så länge innan arbetsgruppen kom samman , med tanke på hur viktig den här frågan är , och vi litade på att den här kommissionen redan från starten skulle börja eftersträva en större jämlikhet mellan kvinnor och män .
jag hoppas att det kommer att ske en förändring och att sammankomsterna blir täta , för det finns många frågor som kommissionen måste ta itu med , så att de åtgärder som leder till en större jämlikhet mellan kvinnor och män påskyndas och leder till goda resultat så snart som möjligt .
fru ledamot , här rör det sig om en uppmaning och inte om en fråga .
men om fru kommissionären vill ge någon förklaring eller visa sin goda vilja ...
låt mig bara få säga en sak till : jag håller med om att kommissionen borde ha sammanträtt tidigare , men förseningen kompenseras av innehållet i sammanträdet , för vi fattade genast viktiga beslut .
fråga nr 39 från ( h-0807 / 99 ) :
angående : gemenskapsinitiativet equal den 13 oktober 1999 antog kommissionen gemenskapsinitiativet equal som syftar till att främja gränsöverskridande samarbete och till att finna och utveckla nya sätt att bekämpa diskriminering och ojämlikhet som på arbetsmarknaden . initiativet är främst inriktat på asylsökande .
inom ramen för detta initiativ skall varje medlemsstat lägga fram förslag i form av ett gemenskapsinitiativ som omfattar den egna staten .
vilka kriterier kommer kommissionen att grunda sig på för att godkänna eller avslå medlemsstaternas föreslagna program ?
vilket gemenskapsorgan skall kontrollera finansieringen av den verkställande kommittén och uppföljningskommittén , och att programmet genomförs på ett riktigt och oklanderligt sätt ?
anslagen från europeiska socialfonden kommer för perioden 2000-2006 totalt att uppgå till 2,487 miljarder euro .
hur mycket kommer grekland själv att bidra med tanke på att gemenskapsinitiativet equal är ett initiativ som förutsätter samfinansiering från medlemsstaternas sida ?
initiativet equqal är inte begränsat till vissa grupper av människor .
det gäller hur man skall motverka diskriminering på arbetsplatserna .
beslutet om detta initiativ fattades i berlin , och då beslutade man att det även skall omfatta de yrkesarbetande bland dem som söker asyl .
jag vill framhålla detta som ett viktigt inslag i detta direktiv .
i varje medlemsstat måste gemenskapsinitiativets program överensstämma med de stadgar som gäller europeiska socialfonden , dvs. equqal följer socialfondens stadgar .
det har presenterats för parlamentet , och vi väntar på parlamentets yttrande i nästa månad .
jag måste betona att initiativet equal svarar mot nationella behov och nationell planering i enlighet med den överenskomna europeiska strategin .
det är i första hand de nationella regeringarna som har ansvaret för att inrätta de gemensamma organen och lägga fram förslag och utse dem som skall genomföra programmen , men det är också i första hand de nationella regeringarna som skall ansvara för kontrollen .
inom europeiska kommissionen finns generaldirektoratet för sysselsättning , som ansvarar för genomförandet , och budgetkontrollen utövas av generaldirektoratet för budgetkontroll , av europeiska byrån för bedrägeribekämpning och av europeiska revisionsrätten .
slutligen har vi frågan om vilken summa som har betalats ut .
grekland har fått 98 miljoner ecu med krav på 80 procents medfinansiering .
för öregionerna och framför allt för de mest avlägset belägna grekiska öarna uppgår initiativets andel till 85 procent och medfinansieringen uppgår till 15 procent .
herr talman ! jag anser att riktlinjerna för gemenskapsinitiativet equal , och speciellt de fyra åtgärder som beskrivs i det , leder till ett mycket komplicerat , byråkratiskt , men egendomligt nog också svåröverskådligt system .
man frågar sig t.ex. på vilket sätt ett utvecklingssamarbete skall bevisa att det är representativt och präglas av samarbetsanda , såsom krävs av åtgärd 2 i artikel 33 i direktiven .
kravet på mellanstatligt samarbete och de komplicerade kraven på planering och genomförande av ett utvecklingssamarbete leder ofrånkomligt tanken till stora system , som ensamma kan uppfylla dessa krav .
detta strider emellertid mot de allmänna målens uttalade önskemål om decentraliserade handlingsplaner , helst på den lokala självstyrelsens eller jordbruksområdenas nivå .
när det gäller de mest utsatta grupperna , såsom asylsökande , invandrare och andra , innebär det att deras medverkan är omöjlig eller bara symbolisk .
om man tänker på att den totala summan är ganska liten - 2,8 miljarder euro för så ambitiösa mål i 15 stater - är jag rädd att det enda vi till sist kommer att kunna bevisa är att arbetslösheten är av ondo .
först skulle jag vilja säga att det skulle vara till stor hjälp för mig , när vi nu behandlar frågan i parlamentet , om ni ville framföra konkreta förslag , som jag kan ta ställning till .
för det andra måste jag säga att initiativet equal varken avser eller kan minska arbetslösheten eller stödja sysselsättningsfrämjande åtgärder .
för detta ändamål finns den europeiska sysselsättningsstrategin och europeiska socialfonden , som förfogar över mycket stora summor och utomordentligt stora resurser , i synnerhet för länder som grekland .
initiativet equal har en konkret uppgift .
att hjälpa till med att få fram statistiskt material , att genomföra undersökningar och inrätta organ som skall kunna stödja de grupper inom befolkningen som drabbats av diskriminering .
vad vi eftersträvar är alltså samarbete mellan lokala grupper , organ för lokal självstyrelse , mellan länder , så att ett erfarenhetsutbyte kommer till stånd . vi vill alltså framför allt att länderna skall utbyta erfarenheter med varandra .
det är dessa tankar som ligger till grund för initiativet och som också avspeglas i dess budget . vårt mål är att samarbetet i största möjliga utsträckning skall omfatta utvecklingsprogram , privata organisationer , lokala myndigheter , för att komma så nära medborgarna som möjligt .
fråga nr 40 från ( h-0808 / 99 ) :
angående : artikel 13 i eu-fördraget och sysselsättning det förslag till kommissionens direktiv som fastställer en allmän ram för likabehandling inom ramen för anställning och sysselsättning , beviljar undantag för religiösa organisationer ( artikel 4.2 ) .
kan kommissionen informera parlamentet om vilka situationer och grupper inom ramen för artikel 13 ( eu-fördraget ) som kan påverkas av ett sådant undantag ?
för en månad sedan lade kommissionen fram ett förslag i frågan om lika behandling i arbetslivet , i överensstämmelse med fördragets uppdrag att genomföra artikel 13 .
förbud mot diskriminering är ledstjärnan i vårt paket med direktiv och program .
men efter förslag från kommissionen och efter ungefär två års överläggningar med arbetsmarknadens parter , med medlemsstaterna , med europaparlamentet , finns det vissa undantag .
och dessa undantag gäller de yrken som måste utövas av personer med en specialiserad yrkesutbildning .
och jag kan ge ett mycket konkret exempel för att förtydliga .
i en religiös skola är det rimligt att man begär och beviljas undantag , med innebörden att den lärare som tjänstgör vid den aktuella skolan skall omfatta samma konfession som skolan .
undantagen är alltså av detta slag .
det rör sig inte om generella undantag , utan dessa skillnader i fråga om behandling i enlighet med de olika medlemsstaternas specialbestämmelser är berättigade endast när det gäller denna specialiserade yrkesutbildning .
detta är en snedvriden tolkning av hur man stoppar diskriminering .
till exempel skulle det vara helt i sin ordning om religiösa skolor sade till en katolik : vi vill inte anställa dig för du är homosexuell .
det vi har här från kommissionen är en förstärkning av en förtryckande hierarki .
det vi borde göra är ju , och jag hoppas ni instämmer herr kommissionär , att anställa människor på grundval av deras kompetens och inte bevara ett sådant bigotteri och en sådan fördomsfullhet , oavsett hur starkt övertygad man än är .
( el ) jag vill betona att detta undantag inte innebär att man kan vägra en person anställning av vilket skäl som helst . av det skäl ni nämnde , på grund av sexuell läggning , etnisk diskriminering eller vad det vara månde .
undantaget ger en möjlighet till urval endast i de fall då det krävs speciell kompetens , som har ett direkt samband med verksamheten .
det är alltså fråga om positiv diskriminering .
i det exempel ni nämnde , i den katolska skolan , är det logiskt att läraren skall vara katolik .
det är bara undantag av detta slag som kan accepteras .
fråga nr 41 från ( h-0813 / 99 ) :
angående : främjande av sysselsättning för kvinnor i starkt missgynnade regioner kvinnor som lever i starkt missgynnade regioner har ofta enorma svårigheter att få arbete . de har i många fall inte något minimikapital och i deras miljö saknas företagaranda , kooperativa traditioner och utbildningsmöjligheter .
vilka åtgärder planeras för att hjälpa dessa kvinnor att överbrygga hinder som hänger samman med deras sociala bakgrund ? har kommissionen för avsikt att lägga fram en politik som säkerställer en miniminivå , för att på ett korrekt sätt återspegla de extrema förhållanden som dessa kvinnor faktiskt lever under , eller kommer deras svåra situation att återigen förbigås i den nya sysselsättningspolitiken ?
för de eftersatta områdena i europa finns ju sammanhållningspolitiken , och för att genomföra denna politik finns samarbetet och de gemensamma insatserna av både strukturfonderna och europeiska socialfonden och jordbruksfonden .
jag vill tala om att de tillgängliga resurserna för problemområdena utgör en tredjedel av den totala budgeten .
dessa regionalpolitiska insatser som utförs enligt gemensamt överenskomna europeiska riktlinjer i varje medlemsstat - dvs. varje medlemsstat har ansvaret för att genomföra detta program - syftar till att öka antalet arbetstillfällen för både män och kvinnor .
jag kan tala om att 70 procent av bidragen för perioden 2000-2006 , som uppgår till 195 miljarder euro , kommer att gå till de mest eftersatta regionerna i europa .
när det nu speciellt gäller kvinnornas möjligheter till förvärvsarbete , vill jag säga , för det första , att socialfonden innehåller en hel pelare med åtgärder som medlemsstaterna måste vidta för att skapa jämställdhet i fråga om arbetstillfällen , dvs. speciella politiska åtgärder som finansieras av socialfonden och gäller kvinnor .
för det andra , i initiativet leader , som just nu är föremål för granskning , prioriterar man särskilt de utvecklingsstrategier som speciellt syftar till att stödja kvinnor i småföretag inom jordbrukssektorn , inom agroturismen , för att sysselsättningen för kvinnor i jordbruksområdena skall öka .
tack fru kommissionär . ni har gett mig ett välment och precist svar i ordalag som jag uppskattar .
ändå kan jag försäkra er om att vi med de medel som finns tillgängliga - och som ni nämner - inte kan nå de missgynnade regionerna .
för det är regioner där bristerna tar överhanden , och de bör likställas med sådana regioner där vi arbetar i ett partnerskap , där det i princip råder brist på allting .
därför undrar jag om ni inte kan undersöka möjligheten att politiken med mikrokrediter , som har gett resultat för partnerskapet , kan tillämpas bland kvinnor i starkt missgynnade regioner , där de har alla odds emot sig .
jag känner väl till de program ni nämner .
jag kan försäkra er om att vi med hjälp av dessa inte når dit där behoven är som störst .
med hjälp av strukturpolitiken - som jag är väl förtrogen med - och med leader och utvecklingen på landsbygden kan vi inte , vilket behövs , främja sysselsättningen bland kvinnor i de missgynnade regionerna .
därför ber jag att ni undersöker möjligheten att en politik med mikrokrediter tillämpas .
kommissionären instämmer och lovat att lägga izquierdo rojos anförande på minnet .
fråga nr 42 från ( h-0817 / 99 ) :
angående : kommissionens planer beträffande presenterandet av ett nytt socialt handlingsprogram det är angeläget att kommissionen snarast presenterar ett nytt socialt handlingsprogram vari en konkret plan redovisas , inklusive tidtabell för genomförande för såväl det lagstiftande arbetet inom området för social trygghet som initiativ till ramavtal inom ramen för den sociala dialogen .
kan kommissionen redogöra för sina konkreta avsikter vad gäller framläggandet av ett nytt socialt handlingsprogram ?
jag räknar med att det nya programmet för kommissionens socialpolitik under nästa femårsperiod kommer att vara färdigt i slutet av sommaren år 2000 .
för att detta program skall bli färdigt och för att vi skall kunna presentera det , bör vi först slutföra överläggningarna med parlamentet , med arbetsmarknadens parter och med de icke-statliga organisationerna .
det är en diskussion som börjar nu , men vi bör ta hänsyn till resultaten från lissabonmötet .
vid europeiska rådets möte i lissabon görs ett nytt försök att ta itu med frågan om den sociala utslagningen , den sociala utslagningens samband med informationssamhället , med den ekonomiska politiken och med reformerna .
dessa resultat kommer att vara mycket viktiga för den slutliga utformningen av kommissionens sociala program .
jag har redan tidigare nämnt för europaparlamentet att ett möte mellan parlamentet och kommissionen kommer att hållas efter lissabonmötet för att diskutera alla aspekter i fråga om den slutliga utformningen av det sociala programmet för perioden 2000-2006 .
det är klart att ett kommande socialt handlingsprogram skall ta hänsyn till utvecklingen , t.ex. inom informationsteknologin , och vara ett modernt socialt handlingsprogram i tiden .
men kan ni också bekräfta det som jag tar upp i min fråga , nämligen att programmet kommer att få en sådan utformning att vi får en konkret tidtabell för de olika typer av lagstiftning på det sociala området , som kommissionen planerar , samt för de initiativ som kommissionen planerar när det gäller den sociala dialogen mellan arbetsmarknadens parter .
vi har ett behov av att se vilka konkreta alternativ kommissionen kommer att ta upp under den kommande perioden och vilka initiativ till avtal den kommer att ta .
jag delar helt er uppfattning , för det första , om att man skall ta hänsyn till informationssamhället - det nämnde jag också .
den sociala utslagningen , kvinnoprogrammet , våra satsningar i fråga om de sociala trygghetssystemen , allt detta måste man nu betrakta ur det nya perspektiv som informationssamhället innebär .
för det andra ; för de initiativ som tas kommer det naturligtvis att finnas en tidsplan för genomförande och systematisk uppföljning .
det finns en punkt där jag inte kan göra några bindande uttalanden , och det gäller lagstiftningen på socialförsäkringsområdet . som ni vet , omfattas denna inte av fördragets artiklar , dvs. fördraget innehåller ingen rättslig grund för socialförsäkringsområdet .
fråga nr 44 från ( h-0819 / 99 ) :
angående : handikappades möjligheter att ta del av den fria rörligheten inom eu i enlighet med artikel 13 amsterdamfördraget skall varje eu-medborgare kunna ta del av den fria rörligheten inom unionen .
för personer med olika slags fysiska handikapp , i behov av särskilda transporter och personlig assistans , är dock denna fria rörlighet fortfarande mycket begränsad .
vilka åtgärder vidtar kommissionen för att underlätta de handikappades möjligheter på detta område ?
den 26 november 1999 godkände europeiska kommissionen ett åtgärdspaket för bekämpning av diskriminering .
när det gäller detta paket och personer med funktionshinder , finns det ett direktiv , som går ut på att bekämpa diskriminering , speciellt på arbetsplatserna .
europeiska kommissionen tror att detta initiativ för bekämpning av diskriminering kommer att bidra till en högre sysselsättningsgrad för personer med funktionshinder och slutligen kommer att underlätta dessa personers fria rörlighet .
det är naturligtvis särskilt viktigt att personer med funktionshinder får tillgång till kommunikationer , myndigheter och alla slags inrättningar , så att personer med funktionshinder får möjlighet till fri rörlighet .
europeiska kommissionen har godkänt ett förslag till direktiv om specialbestämmelser för bussar , långfärdsbussar och andra fordon , så att dessa blir tillgängliga även för rörelsehindrade personer , inklusive rullstolsburna .
dessutom kan jag meddela att rådet den 4 juni 1998 godkände en rekommendation om att införa en typ av alleuropeiskt parkeringskort för personer med funktionshinder , och syftet med rekommendationen är att hjälpa dem att röra sig fritt i alla medlemsländerna med hjälp av ett gemensamt parkeringskort , så att de kan utnyttja alla anordnade parkeringsplatser i europa .
min fråga rör i första hand handikappades möjligheter att passera gränserna i europa .
det är en ganska dyr historia om man skall ta sig från göteborg till någon plats i övriga europa på semester eller på studiebesök om man sitter i rullstol och dessutom behöver ha med sig en personlig assistent eller medhjälpare för att klara av situationen .
jag är tacksam över att kommissionen har antagit en handlingsplan .
det är ju emellertid en förutsättning att det finns ekonomiska resurser och möjligheter att rent fysiskt komma över gränserna om man har ett funktionshinder .
det skulle vara intressant att höra om kommissionen också är beredd att avsätta ekonomiska medel för de personer som har funktionshinder , så att också de skall kunna ta sig längre ut i världen än dit rullstolen tar dem .
jag nämnde kommissionens förslag till direktiv om att de allmänna kommunikationerna måste utformas så att de kan utnyttjas av personer med funktionshinder .
rådet har inte tagit ställning till förslaget , som är föremål för överläggningar .
jag anser att ett sådant strategiskt beslut kan fattas på europeisk nivå .
det är enligt min mening utomordentligt svårt med en specialinriktning för att lösa varje enskild persons transportproblem .
detta oavsett om det gäller specialprogrammen för utbildning , för ungdomar och kvinnor eller om det måste genomföras genom nationell politik .
fråga nr 45 från ( h-0006 / 00 ) :
angående : genomförande av direktiv 96 / 71 / eg om utstationering av arbetstagare direktivet om utstationering har ännu inte genomförts i danmark trots att tidsfristen har löpt ut .
det lagförslag som lagts fram i folketinget innehåller inga bestämmelser som reglerar lönearbetsrättigheter enligt kollektivavtal .
enligt artikel 3.8 i direktivet skall arbets- och anställningsvillkor vara i överensstämmelse med de &quot; kollektivavtal som har ingåtts av de mest representativa arbetsmarknadsorganisationerna på nationell nivå och som gäller inom hela det nationella territoriet &quot; .
en sådan användning av ett avtal utanför dess individuella område kan emellertid inte åläggas parterna utan stöd i lagen .
det finns därför två möjliga lösningar : antingen gäller direktivet inte i danmark eller så innebär direktivet att danmark måste införa allmängiltiga avtal .
kan kommissionen bekräfta att direktivet om utstationering inte gäller i danmark beträffande &quot; kollektivavtal &quot; med &quot; allmän giltighet &quot; ( se artikel 3.1 ) eftersom sådana avtal med allmän giltighet inte existerar i dansk rätt ?
om inte , hur skall direktivet uppfyllas på denna punkt ?
europeiska unionens direktiv om utlandsplacering av arbetstagare innebär att samma arbetsvillkor som gäller för mottagarlandet också skall gälla för de utländska arbetstagare som placerats i detta land .
direktivet innebär att två regelsystem kan tillämpas : antingen mottagarlandets lagstiftning eller de kollektivavtal som tillämpas generellt inom en viss bransch .
eftersom danmark inte har ett system som innebär att kollektivavtal upphöjs till allmänt gällande regler , måste man vid tillämpningen av lagstiftningen räkna med att inte bara lagstiftningen om arbetsvillkor utan också de allmänt tillämpliga kollektivavtal som slutits av de mest representativa organisationerna gäller för de utlandsplacerade arbetstagarna .
enkelt uttryckt kan man alltså säga att danmark har två alternativ ; antingen att stifta lagar eller också att välja ut ett kollektivavtal och ge det status av lag .
det förs en diskussion mellan europeiska kommissionen och danmark , och vi räknar med att danmark skall meddela när detta direktiv har införlivats i dess nationella lagstiftning .
danmarks tidsfrist för att besvara kommissionens frågor löpte ut den 6 december 1999 . vi har inte fått något svar .
vi avvaktar för att se vilka steg som kommer att tas i fortsättningen .
tack för ett mycket tydligt svar som - om tolkningen stämmer - innebär att direktivet om utstationering medför en skyldighet för danska staten att inrätta ett system med allmänt användbara avtal .
det är ett mycket tydligt svar , men det är också ett svar - vilket jag måste göra er uppmärksam på - som ställer de danska organisationerna , den danska regeringen och det danska folketinget i en politiskt sett mycket , mycket svår situation , eftersom det är känt att det finns några grundläggande problem i förhållandet mellan den danska modellen som i hög grad bygger på kollektiva avtal , och den kontinentala modellen som förutsätter lagstiftning .
den oenighet och korrespondens som ni , fru kommissionsledamot , hänvisar till , rör ju först och främst ett annat direktiv , dvs. arbetstidsdirektivet , men nu kan vi alltså se fram emot en ny uppmaningsskrivelse och kommande domstolsförhandlingar som ett resultat av att den danska regeringen inte kommer att , eller uttryckligen har meddelat , att man inte har för avsikt att genomföra lagstiftning och tillämpa allmänt användbara avtal .
för det första ; vi försöker inte ändra systemet vare sig i danmark eller i något annat land .
som jag svarade tidigare , finns det alltid problem när det gäller tolkningen av europeiska kommissionens direktiv , dels därför att de är mycket allmänt hållna , men dels också därför att systemen skiljer sig mycket mellan de olika länderna .
när det gäller er fråga , kan jag säga att det konkreta problemet inte bara gäller danmark .
det är inte bara danmark som har olösta frågor .
fem länder har införlivat direktivet i sin nationella lagstiftning , och i de övriga pågår diskussioner .
det har förts diskussioner mellan kommissionen och den danska regeringen men också de andra regeringarna , därför att man måste hitta den bästa metoden för att utlandsplacerade arbetstagare i danmark skall omfattas av beslut som fattats på europeisk nivå av alla medlemsländerna .
vi räknar med att både danmarks och ytterligare nio länders regeringar skall vidta åtgärder i denna riktning .
tack fru kommissionär för det engagemang ni har visat .
ni har lyckats uppnå dagens mål : att besvara samtliga frågar .
eftersom tiden för frågestunden med frågor till kommissionen är över , kommer frågorna nr 46 och 68 att besvaras skriftligen .
ansvarsfrihet 1997
nästa punkt på föredragningslistan är betänkande ( a5-0004 / 2000 ) av van der laan för budgetkontrollutskottet om beviljande av ansvarsfrihet för kommissionen och om avslutningen av räkenskaperna för europeiska gemenskapernas allmänna budget för budgetåret 1997 ( avsnitten i - parlamentet , ii - rådet , iii - kommissionen , iv - domstolen , v - revisionsrätten ) ( sek ( 1998 ) 520 - c4-0350 / 1998 , sek ( 1998 ) 522 - c4-0351 / 1998 , sek ( 1998 ) 519 - c4-0352 / 1999 ) .
kommissionären är ännu inte här , men jag hoppas och antar att hon kommer om ett par minuter .
jag vill föreslå att vi börjar trots detta , och hoppas att kommissionären , om hon fortfarande är kvar på sitt kontor , kan lyssna till talet , i synnerhet föredragandens tal .
herr talman ! fru schreyer har säkerligen ett mycket gott skäl för att inte vara här , för annars skulle hennes frånvaro vara oförlåtlig .
jag skulle vilja börja med att tacka mina kolleger för deras medverkan till detta betänkande . det skulle inte ha varit vad det är i dag utan denna samarbetsanda .
herr talman ! i början av förra året sköts beviljandet av ansvarsfriheten för 1997 upp , eftersom parlamentet omöjligen kunde bevilja ansvarsfrihet åt en avgående kommission som inte skulle kunna åta sig förpliktelser för framtiden .
i sin resolution hävdade parlamentet att ansvarsfrihet skulle kunna beviljas först efter det att vi fått seriösa , långtgående reformförslag från den nya europeiska kommissionen .
detta betänkande läggs nu fram vid en avgörande tidpunkt , omedelbart före kinnocks reformer .
det är en utmärkt chans för parlamentet att sätta en långtgående reformstämpel på dessa planer .
redan under förarbetet har det visat sig att kommissionen på grundval av de första utkasten kommit med mycket viktiga löften .
vi krävde en föreskrift för &quot; angivare &quot; , och en sådan har kommit .
parlamentet ville ha en åtskillnad mellan ekonomistyrning och revisionsfunktioner .
den har vi redan uppnått .
parlamentet kräver en uppförandekod för kommissionärer och kabinett .
även det har vi fått .
parlamentet bad kommissionen att avstå från sina överdrivna förmåner .
även detta har de gjort .
samtidigt har kommissionen förpliktigat sig att samarbeta med parlamentet på området sem-2000 .
man kommer också att se över kontoren för tekniskt bistånd för att vidta grundläggande förändringar .
detta är några goda första steg som visar att , om parlamentet så vill , förändringar inte bara är möjliga utan också snabbt kan omsättas i handling .
vi vill dock ännu mer .
kommissionen måste nu komma med ett ambitiöst och långtgående reformprogram .
det är inte bara nödvändigt för en oklanderlig offentlig förvaltning ; det är en conditio sine qua non för att återställa förtroendet hos medborgarna i europa .
vi kräver nu tydliga löften av europeiska kommissionen på följande punkter .
för det första måste parlamentet få fullständig tillgång till kommissionens samtliga handlingar .
detta står visserligen i motsats till att vi internt snabbt måste nå en uppgörelse för att kunna garantera sekretessen för känsliga dokument .
i samband med inhämtande av information skulle jag vilja göra kommissionen uppmärksam på att vi är mycket oroliga över de preliminära planer som föreligger om allmänhetens tillgång till handlingar .
om det aktuella utkastet kommer att gå igenom är det ett oerhört steg tillbaka jämfört med i dag .
det måste bli slut på en situation där finansiellt starka organisationer med representanter i bryssel kan komma åt information men inte de vanliga medborgarna .
det får inte heller vara så att en offentlig institution innehar copyright till offentliga handlingar .
vidare vill vi ha tydliga arbetsbeskrivningar för varje europatjänsteman så att en tjänsteman har dessa samvetsskäl och lättare kan opponera sig mot uppdrag som är oetiska eller olagliga .
vidare måste det vara så att när revisionsrätten upptäcker att en brist uppträder inte bara ett år utan två år efter varandra bär förvaltningen ansvar för detta , och sådant skall även kunna gå ut över en karriärplanering .
slutligen måste vi naturligtvis också ha ett bättre samarbete mellan europeiska revisionsrätten och dess nationella motparter .
parlamentet kräver också av kommissionen att den den 31 mars i år kommer med en första skiss för reformeringen av den externa biståndspolitiken .
det får inte längre vara så att europa visserligen är en ekonomisk makt men att vi inte har något politiskt inflytande därför att vi , när det kommer till kritan , inte kan erbjuda någon effektiv hjälp till områden som verkligen är i behov av sådan .
som exempel på detta nämner jag gaza .
det är oacceptabelt att kommissionen färdigställde ett sjukhus 1996 och att det ända fram till den dag som i dag är inte har legat en enda patient i det .
herr talman ! sedan 1996 har ansvarsfriheten fått en tung politisk betydelse .
det är ett av de starkaste maktmedlen som parlamentet har , och därför måste det användas med försiktighet .
därför kommer vi med all sannolikhet att bevilja ansvarsfrihet i morgon .
vi avhänder oss dock inte detta vapen utan att också placera ut en tidsinställd bomb .
ansvarsfriheten för 1999 kommer nämligen att beviljas först när alla de ekonomiska oegentligheter som revisionsrätten upptäckt har lösts .
slutligen , denna ansvarsfrihetsrapport riktar sig naturligtvis också till kommissionen .
men det hindrar inte att också europaparlamentet måste får ordning på torpet internt .
så länge vi inte har någon stadga är vi inte trovärdiga som unionens reformeringsmotor .
reformerna av de europeiska institutionerna är ett nödvändigt villkor för att kunna bygga vidare på europa .
det enda sättet att få ett handlingskraftigt och rättvist europa är att också se till att det är öppet och demokratiskt .
alla institutioner måste nu slå sig ihop för att tillsammans arbeta för ett sådant europa .
( en ) herr talman ! utskottet för industrifrågor bestämde sig för att upprätta ett betänkande om ansvarsfrihet för 1997 trots att vi inte särskilt har ombetts att göra det .
vi gjorde detta eftersom vi tyckte att vi borde inleda denna mandatperiod på det sätt vi har för avsikt att fortsätta den , det vill säga genom att se till att vi tar väl hand om skattebetalarnas pengar i europa .
under vårt arbete på detta betänkande stod det klart att det finns kvarhängande problem inom de utgiftssektorer som ligger i vår budget .
de är inte unika för 1997 och verkar ha två röda trådar .
den första är kommissionens tendens att ge sig in på mycket ambitiösa program , särskilt i tredje världen , utan att tillräckligt ha utvärderat de praktiska detaljerna kring genomförandet och utan ordentlig resurstilldelning .
den andra gäller allvarliga administrativa brister hos kommissionen , särskilt vad beträffar samordningen mellan avdelningar och hanteringen av externa kontakter .
jag vet att alla institutioner har del i ansvaret för kommissionens ökade arbetsbörda och för en del av resursbristen .
det kan inte ursäkta allt det vi har stött på .
europas medborgare förväntar sig att de europeiska institutionerna administreras ordentligt och det gör de rätt i .
det är därför jag vill upprepa min kollegas kommentarer om vikten av den reformprocess som herrar prodi och kinnock har lovat europas folk .
att döma av det jag har sett av reformprocessen ser det bra ut .
jag såg några av kinnocks papper i dag och jag hörde en del av det han hade att säga .
jag är full av tillförsikt om att vi och europas politiker kommer att få den slags reform vi behöver om vi stöder honom .
men vi behöver denna reformprocess .
många av de generella punkter som tas upp i vårt utskotts betänkande omfattas av van der laans betänkande .
det är ett utmärkt betänkande och vi bör alla gratulera henne till det .
jag tycker att man verkar ha hittat alla de ömma punkterna utan att betänkandet bara blir en uppsättning detaljer , som några av de gamla betänkandena .
de grupperas samman och detta är mycket viktigt .
jag skulle vilja fästa er uppmärksamhet på två frågor .
den ena är kärnkraftssäkerhet i östeuropa .
vi måste få ordning på detta .
den oberoende expertkommittén sade att kommissionen inte skötte detta ordentligt .
vi måste råda bot på detta .
den andra punkten gäller granskningsmekanismer .
vi behöver ha material från kommissionen som vi kan använda som hjälp vid granskningen av utgifterna .
vi behöver ordentlig information som lämnas på rätt sätt och vi måste alla ta hela denna process mycket mer på allvar än vi har gjort hittills .
den har betraktats som en byråkratisk process som skulle göras så snabbt som möjligt med så liten tidsåtgång som möjligt .
jag hoppas att kollegerna i denna kammare kommer att stödja skälen för ansvarsfrihet för 1997 och att samtidigt kommissionen kommer att driva på reformprocessen som borde ha genomförts för länge sedan .
det är enda sättet att skapa en ny kultur i kommissionen och samtidigt återställa allmänhetens förtroende .
herr talman ! jag är säker på att kommissionen kommer att bli lättad över att höra att ansvarsfriheten för 1997 troligen inte kommer att få samma konsekvenser som ansvarsfriheten för 1996 vilken , som ni alla är så väl medvetna om , ledde till att santer-kommissionen tvingades avgå .
socialistgruppen kommer att rösta för ansvarsfrihet .
jag är säker på att ni blir lättade av att höra också detta .
men därmed inte sagt att vi är nöjda , därmed inte sagt att allt är rosenrött .
det står klart att en radikal omvälvning av kommissionen borde ha gjorts för länge sedan .
detta betyder emellertid att vi erkänner att de åtgärder man vidtar går i rätt riktning .
jag vill bara skissera några av de frågor där vi socialister har föreslagit ändringar .
vi hoppas att dessa kommer att bifallas eftersom de är viktiga på grund av sin inverkan på den kommande reformen .
för det första tjänstemännens immunitet : denna bör upphävas om och när en nationell åklagare så begär .
vi måste göra det mycket lättare att åtala tjänstemän som har gjort sig skyldiga till bedrägeri och korruption .
det är avgörande att man noterar att kommissionen allt för ofta har underlåtit att genomföra de reformer som revisionsrätten har rekommenderat .
det finns skäl till att rättens rapport finns , det finns skäl till vårt svar och det är viktigt att det följs upp .
jag hörde just att kommissionen kommer att inrätta en arbetsgrupp för revisionsuppföljning .
så även om vi inte hör någonting mer vet vi att det går åt rätt håll vad beträffar de reformer vi vill ha .
allt för ofta har vi lagt fram rekommendationer och de har inte lett till någon åtgärd , trots att ni väldigt ofta har sagt att ni skulle handla i enlighet med dem .
vi vill se denna uppföljning i mycket större utsträckning i framtiden .
den andra frågan är tillgången till konfidentiella handlingar .
vi har tidigare haft problem i fråga om vår skyldighet att ta ställning till ansvarsfrihet eftersom vi inte har haft tillgång till de handlingar vi borde ha haft .
vi inser att även vi har ett ansvar här , att om vi får handlingar måste vi tillse att sekretessbelagda handlingar verkligen förblir sekretessbelagda .
en fråga som man hänvisar till i van der laans betänkande är hela frågan om sjukhuset i gaza .
situationen där är helt oacceptabel .
vi kommer inte att tolerera den mycket längre och vi vill att man omedelbart agerar i denna fråga .
jag skulle vilja gratulera lousewies van der laan .
vanligtvis bryr jag mig inte om att gratulera människor , men jag tycker att hon har producerat ett mycket övertygande betänkande och förtjänar vårt tack .
herr talman , kolleger , fru kommissionär ! låt oss vara ärliga ; vi befinner oss i en något märklig situation .
vi diskuterar ansvarsfrihet för ett år som ligger bakom oss , men vi diskuterar också kommissionens ansvar .
jag vill ta upp de problem som fortfarande ligger i skyhöga travar på vårt bord .
bedömningen i fråga om att bevilja ansvarsfrihet eller inte hänger också i viss mån samman med var man lägger den största tonvikten .
det handlar om en kommission som inte längre sitter kvar .
det är en ny kommission .
då är det logiskt att bevilja ansvarsfrihet , för vad kan den nuvarande kommissionären förebrås för när det handlar om året 1997 ?
de problem som är aktuella finns fortfarande kvar , och då börjar man att tvivla .
vi måste nu fatta ett beslut om kommissionens goda föresatser , men det föreligger fortfarande ingen strukturerad översikt över dessa goda föresatser .
kinnock kommer med sitt förslag nästa månad .
det väntar vi allesammans med spänning på , men vi har ännu inte den kunskapen när vi nu måste fatta beslut om ansvarsfrihet .
det är tydligen ett dilemma som föredraganden också har brottats med .
detta dilemma är ännu mer vidsträckt än de områden som jag nämnde .
det handlar till exempel om kommissionens löften .
de ser i sig bra ut .
jag har läst ett antal av kinnocks dokument , och de har vi fullt förtroende för .
men jag ger två exempel på varför det inte är självklart att de goda föresatser som kommissionen nu gett uttryck för kommer att leda till ett gott resultat . offentligheten , sekretessbelagda handlingar .
detta togs också upp av föregående talare .
det cirkulerar nu ett dokument , inte på låg nivå utan på hög nivå i kommissionen , varvid offentligheten för dokument inte utökas utan helt enkelt upphävs .
ett exempel på att ett vackert löfte inte automatiskt kommer att leda till ett gott resultat .
det gäller också för &quot; angivarna &quot; .
kinnock har också ägnat dem några vackra ord , men samtidigt är det fullständigt otydligt , just nu när vi skall fatta beslut om detta , vad som till exempel händer med &quot; angivare &quot; som inte får någon chans internt utan som vill gå ut , till pressen , till parlamentet .
det har fortfarande inte kommit något svar på den sortens avgörande frågor på det området .
det råder således tvivel , just nu när vi skall fatta beslut om detta , om dessa löften från kommissionen är tillräckligt kraftfulla .
detta gäller också till exempel för de mycket konkreta projekt som utskottet för industrifrågor har tagit upp .
jag anser att kommissionen och kinnock måste komma med goda föresatser , med goda planer för personalpolitiken , för den ekonomiska förvaltningen , men varje kommissionär som nu är ansvarig för ett område med allvarliga brister i det förflutna måste komma med goda planer för att förbättra situationen och inte med allmänna vackra förslag .
för närvarande har vår grupp fortfarande förbarmande , tålamod med kommissionen eftersom den inte kan ställas till ansvar för många felaktigheter ur det förflutna , men detta tålamod är inte obegränsat .
det måste finnas tydliga framsteg i sikte .
för närvarande förlitar vi oss på att kommissionen kommer med dessa goda förslag , men detta förtroende är inte automatiskt .
slutligen , herr talman , ansvarsfriheten 1996 var början till slutet för den förra kommissionen .
jag uttalar förhoppningen , men ännu starkare , jag vill egentligen kräva av den nuvarande kommissionen att ansvarsbefrielsen 1997 är inledningen till en verklig reformering av den ekonomiska politiken från kommissionens sida , för annars kommer denna ansvarsbefrielse inte att ha varit till någon nytta .
när man bedömer frågan om ansvarsfrihet för kommissionen , måste avgörandet grundas på vad som faktiskt hände under det aktuella budgetåret , i detta fall under år 1997 .
i vår grupp har vi svårt att se att den ekonomiska förvaltningen för år 1997 på något avgörande sätt var bättre än den för år 1996 .
det året röstade vi mot ansvarsfrihet .
i konsekvens med detta kommer vi att rösta mot ansvarsfrihet även för år 1997 .
vi menar att denna vår bild bekräftas av revisionsrättens granskning .
det är både bra och nödvändigt att reformer har utlovats .
ännu så länge återstår det dock att infria de löften som givits , inte minst vad gäller öppenhet .
vi kommer därför att rösta för de krav på reformer som framförs i resolutionen , men mot att ansvarsfrihet beviljas .
herr talman ! för det första har jag bara positiva ord att säga om van der laans mycket väl utförda arbete i samband med detta betänkande .
gruppen unionen för nationernas europa kan inte rösta för ett godkännande av räkenskaperna för budgetåret 1997 .
betänkandet om s.k. ansvarsfrihet innehåller en omfattande och ytterst kritisk genomgång av räkenskaperna .
vi stöder dessa kritiska anmärkningar och därför måste jag konstatera att det verkar helt absurt mot denna bakgrund att acceptera ett godkännande .
det har inte varit möjligt för revisionsrätten att avge en revisionsförklaring om att de dispositioner som räkenskaperna omfattar är lagliga , och vi anser det vara ytterst problematiskt att vi som ledamöter av detta parlament skulle rösta för räkenskaperna utan att säkert veta om dispositionerna är lagliga .
majoriteten har beviljat ansvarsfrihet under förutsättning att den nya kommissionen genomför en rad reformer som skall se till att det vi erfarit under den förra kommissionens mandatperiod inte upprepas .
jag måste återigen säga att det handlar om en högst olycklig sammanblandning av den gamla kommissionens ansvar för budgetåret 1997 och den nya kommissionens ansvar för framtiden .
vi menar inte att den nya kommissionen under några omständigheter skall ha ansvar för den gamla kommissionens politik .
vi menar att det är felaktigt att tala om kommissionens ansvar som en institution .
bristerna fram till 1999 skall skyllas på de som då hade ansvaret och vi har ännu inte möjlighet att se om den nya kommissionen kan göra det bättre .
i och med detta märkliga förfarande tar inte parlamentet chansen att placera ansvaret för dispositionerna under budgetåret 1997 där det hör hemma , dvs. hos den tidigare kommissionen .
det var 1996 års budget som fällde den tidigare kommissionen och 1997 års budget är precis lika betungande .
det finns inget skäl till att vi mot denna bakgrund skulle bevilja ansvarsfrihet .
vad gäller beslutet om avslutningen av räkenskaperna vill vi inte delta i omröstningen och slutligen vad gäller resolutionsförslaget vill vi betona de många korrekta godkännandena och rösta för .
herr talman ! beslutet om ansvarsfrihet för budgetåret 1997 har skjutits upp , eftersom den kommission som beslutet vid den tidpunkten gällde hade trätt tillbaka och bara var en expeditionskommission .
i dag föreslås det nu i van der laans betänkande - som hon har lagt ned mycken flit på , och det bör man tacka henne hjärtligt för - att kommissionen medges ansvarsfrihet för budgetåret 1997 .
man kan fråga sig varför den nuvarande kommissionen får ansvarsfrihet för hur den förra kommissionens skött sin ekonomi - camre har just berört detta - framför allt som den förvägrades ansvarsfrihet för år 1996 .
men så ligger det till .
i och med att den nya kommissionen övertog mandatet är den också ansvarig för både goda och dåliga prestationer i det förflutna .
eftersom kommissionen till sitt system är ett kollegium och endast kan medges ansvarsfrihet i sin helhet , respektive kan få den uppskjuten eller förvägrad , spelar det inte heller längre någon roll att fyra förutvarande kommissionärer hörde till den tidigare kommissionen som hittills inte medgivits ansvarsfrihet , och nu åter är ledamöter i denna institution .
denna fråga skulle ha behövt ställas när den nya kommissionen tillsattes .
om parlamentet denna vecka röstar för budgetkontrollutskottets förslag och beviljar ansvarsfrihet , får kommissionen inte förstå detta som en check in blanko .
ty enligt min åsikt är den tredje delen i van der laans betänkande den viktigaste , nämligen resolutionsförslaget .
de villkor som samlats under åtta rubriker är väsentliga beståndsdelar av ansvarsfriheten , och vårt beslut utgår från att de uppfylls .
under processen med beviljande av ansvarsfrihet för åren därefter - 1998 är redan påbörjat - kommer parlamentet att mycket noga få lov att undersöka om det inte alltför snabbt gett kommissionen ett förtroendeförskott för år 1997 .
det kommer genast att visa sig , när kommissionen lägger fram sitt reformprogram .
huruvida det då finns någon effektivitet , öppenhet och ansvar , liksom en uttalad informationsvilja gentemot den myndighet som beviljar ansvarsfrihet , kommer vi att granska när ansvarsfrihet för budgetåret 1998 skall beviljas .
herr talman ! vi minns alla att parlamentet beslöt att skjuta upp ansvarsfriheten för budgetåret 1997 i avvaktan på åtaganden från den nya europeiska kommissionen om interna reformer .
som svar på detta har kommissionen gjort olika åtaganden och har helt klart fattat många beslut om reformer .
i rättvisans namn måste man säga att den nye ordföranden prodi och hans lag verkligen har förbundit sig att genomföra de mekanismer för ekonomisk kontroll detta parlament har lagt fram .
reformeringen av europeiska kommissionen måste dock nu ses mot bakgrund av den debatt som kommer att äga rum inför den kommande regeringskonferensen och reformeringen av olika politiska områden och initiativ inom eu .
dagens eu-fördrag kommer att ändras för att till exempel säkerställa att utvidgningen kan lyckas .
jag tvivlar inte på att ytterligare reformer av eu : s institutioner kommer att analyseras i denna debatt .
men ur de små medlemsstaternas perspektiv är det viktigt att europeiska kommissionen reformeras på ett sätt som säkerställer att små medlemsstater fortfarande är företrädda i kommissionen .
herr talman ! nu får kommissionen sin ansvarsfrihet för budgetåret 1997 , men i realiteten förtjänar de den inte .
år 1997 lyder under den gamla kommissionen och därför menar den nya att den inte kan ta på sig ansvaret .
det är korrekt att genomförandet av budgeten för år 1997 härrör till den gamla kommissionen , men den nya kommissionen har i gengäld åtagit sig att rensa upp efter de gamla skandalerna och jag måste erkänna att jag inte är särskilt imponerad .
mentaliteten från förr då man skulle sopa allt under mattan och ställa upp för sina vänner , existerar tyvärr alltjämt .
det finns vissa som menar att vi är bättre betjänta av att begrava gamla synder och börja på ny kula .
jag anser att vi inte kan börja på ny kula om vi inte först rensar upp ordentligt .
jag avser här i synnerhet de gamla skandalerna i echo .
det gör mig mycket irriterad att det är så svårt att få ut handlingar om frågan .
jag är föredragande för echo i budgetkontrollutskottet och det kommer att bli mycket svårt för mig att utföra mitt arbete om inte kommissionen ger mig den nödvändiga informationen .
utifrån ser det ut som om kommissionen har något att dölja .
mina undersökningar tyder dessvärre också på att så skulle kunna vara fallet .
kommissionen lägger inte alla kort på bordet och återupptar alltså sin hävdvunna praxis .
det var denna praxis som ledde fram till kommissionens fall .
jag kan därför fullständigt stödja uppmaningen att parlamentet skall ha tillgång till alla handlingar .
i annat fall kan vi inte utföra vårt arbete .
åtgärder att vidta med anledning av den oberoende expertkommitténs andra rapport
nästa punkt på föredragningslistan är betänkande ( a5-0001 / 2000 ) av van hulten för budgetkontrollutskottet om åtgärder att vidta med anledning av den oberoende expertkommitténs andra rapport om reformering av kommissionen .
( en ) herr talman ! vid den här tiden förra året inrättade europaparlamentet en oberoende expertkommitté med middelhoek som ordförande , som skulle granska anklagelser om bedrägeri , nepotism och korruption i europeiska kommissionen .
15 mars offentliggjorde kommittén sin första rapport med slutsatsen att : &quot; det börjar bli svårt att hitta någon som har någon som helst ansvarskänsla &quot; .
bara några timmar efter det att rapporten hade framlagts tillkännagav ordförande santer att hela hans kollegium avgick .
avgången markerade slutet på en bitter kamp mellan ett allt mer självsäkert parlament och en kommission som var befläckad av skandalanklagelserna .
sedan dess har situationen i bryssel förändrats till oigenkännelighet . ett nytt parlament med en ny vigör har valts och en ny kommission tillsatts .
när den nominerade ordföranden prodi talade i denna kammare 21 juli förband han sig att beakta den andra rapporten från den oberoende expertkommittén för reformering av kommissionen fullt ut . denna innehåller 90 detaljerade rekommendationer och det är den vi diskuterar i dag .
den nya kommissionen har redan tagit viktiga steg bort från sitt gamla sätt att fungera .
en uppförandekod för kommissionärer och deras kabinett har antagits .
som en symbolisk men betydelsefull gest har kommissionärerna frivilligt avstått från sin rätt till skattefria inköp av alkohol , tobak , bensin och konsumentvaror .
nya regler har tagits fram och förverkligats vad beträffar hur högre tjänstemän utses .
antalet avdelningar har minskats .
enligt min mening har kommissionen visat ett tydligt engagemang utan tidigare motstycke för förändring och detta skall de ha en eloge för .
det övergripande syftet med reformerna måste vara att skapa en stark , ärlig europeisk offentlig sektor som är rustad för att genomföra sina uppgifter på ett effektivt och kompetent sätt , en offentlig sektor där tjänstemännen har medel att genomföra sina uppgifter och hålls fullt ansvariga på alla nivåer , en offentlig sektor som känner igen och belönar det förtjänstfulla och uppmuntrar tjänstemännen att utveckla hela sin potential .
för att uppnå detta måste vi agera på fyra områden .
för det första måste den ekonomiska hanteringen och kontrollen inom kommissionen förbättras .
ett av de största problemen är att det saknas ett fungerande system för ekonomisk kontroll .
kommissionens generaldirektorat måste få ett totalansvar för sina egna kostnader , inklusive den ekonomiska kontrollen .
ett nytt oberoende revisionssystem måste införas .
generaldirektoraten måste offentliggöra sina egna årsberättelser så att problemområden tydligt kan identifieras och uppställa årliga mål för att minska bedrägerier och regelbrott .
i utbyte för denna större självständighet måste cheferna göras fullt och personligen ansvariga för sitt agerande .
det är klart att övergången till ett sådant nytt system kommer att ta tid .
det kommer att krävas förändringar i budgetförordningen och parlamentet måste uttala sig om dessa förändringar .
men även om kommissionen måste se till att den följer fördraget och budgetförordningen under en övergångsperiod får inte detta bli en ursäkt för att inte göra någonting .
det finns ett trängande behov av förändringar i dag .
för det andra måste kampen mot bedrägeri , misskötsel och nepotism intensifieras , främst genom att man skapar en kultur där de inte kan frodas .
detta kräver att kommissionärerna och de högre tjänstemännen statuerar klara exempel och erbjuder lämplig utbildning , och dessutom att de befintliga mekanismerna för att hantera bedrägerier förstärks .
olaf , kommissionens byrå som skapades tidigare i år , måste sättas under en oberoende europeisk allmän åklagares ledning , vars uppgift skall vara att förbereda åtal i nationella brottmålsdomstolar av kriminella handlingar som begåtts mot unionens ekonomiska intressen av ledamöter och tjänstemän i de europeiska institutionerna .
ett förslag kan läggas , ett förslag bör läggas , på grundval av artikel 280 i fördraget senast vid halvårsskiftet .
för det tredje måste det europeiska offentliga livet uppfylla högt satta normer .
den politiska kris som ledde till att kommissionen föll tidigare i år visade tydligt på behovet av otvetydiga uppföranderegler vars efterlevnad kan framtvingas .
ett antal koder har sedan införts .
de måste utvärderas av parlamentet och bör göras juridiskt bindande .
de europeiska institutionerna bör följa det exempel som ett antal länder har satt , i synnerhet storbritannien , och tillsätta en kommitté för normer i det offentliga livet med mandat att ge råd om yrkesetik och uppföranderegler inom de europeiska institutionerna .
uppgiftslämnare som är i god tro måste skyddas .
i slutet av förra året tillkännagav kinnock nya åtgärder för att skydda uppgiftslämnare .
dessa måste genomföras utan dröjsmål .
även om sådana åtgärder aldrig kan bli ett alternativ till en god ledning måste det finnas en säkerhetsventil när någonting går fel .
det är avgörande att reformerna inte begränsas till kommissionen .
även parlamentet måste överväga behovet att förbättra sina interna regler , administrativa rutiner och ledningsutövning .
slutligen måste kommissionens personalpolitik moderniseras .
den är helt klart inte anpassad till kraven från en modern , multinationell organisation .
den sociala dialogen har ofta fungerat som en broms för reformer och borde ha setts över för länge sedan .
det måste bli mer attraktivt att arbeta inom de europeiska institutionerna .
allt för många unga , nya tjänstemän lämnar sina jobb efter bara några år .
förtjänster måste erkännas och belönas , specialutbildning måste bli ett sine qua non för befordran till högre befattningar .
befordringssystemet måste göras rättvisare och ges ökad insyn .
sist men inte minst måste löne- och förmånspaketet ses över .
det måste bli flexiblare och visa större ansvar för arbetsmarknadens villkor .
det måste befrias från vissa av sina mest förlegade beståndsdelar och man måste ta itu med den berättigade kritiken från allmänheten , som inte kan inse varför eu : s tjänstemän skall få utflyttningsbidrag i all oändlighet i ett europa med öppna gränser eller betala skatter vars nivå ofta ligger långt under nivån i medlemsstaterna .
kommissionär kinnock kommer att framlägga sitt meddelande om reformerna i morgon .
detta meddelande måste innehålla en klar tidtabell .
med en ny kommission och ett nytt parlament i full gång är incitamentet för reformer starkare än det någonsin har varit och förmodligen någonsin kommer att bli .
utvidgningen av unionen ligger bara några år framåt i tiden .
nu är det dags för europa att göra rent hus och inpränta en ansvarskänsla - som de oberoende experterna kunde ha sagt - hos sina institutioner .
i juni förra året gav väljarna i europa en tydlig signal om att de är trötta på ändlösa historier om misskötsel och nepotism .
det finns ett mycket enkelt sätt att handskas med dessa historier .
låt oss avskaffa misskötsel och nepotism .
herr talman ! jag hoppas verkligen att ingen missförstår mig och därför vill jag först av allt säga att jag naturligtvis är för en kamp mot bedrägeriet och att jag med kraft stöder alla lämpliga och nödvändiga reformer .
detta är en fråga som inte är enkel och som skulle behöva fördjupas betydligt mer , men jag kommer att nöja mig med att bara peka på enstaka punkter , bl.a. för att ni , om möjligt , skall bli medvetna om vad vi talar om .
experterna kan ge information och upplysningar , formulera uppfattningar och ge råd , men de har inte något politiskt ansvar gentemot sina väljare .
i stället är det politikerna som måste undersöka vad de kan utnyttja i en expertrapport och vad man inte kan tillämpa i sin helhet i en anda av , som det ibland har verkat , självplågeri .
jag tror - låt mig bara nämna ett par punkter - att när det gäller ledamöterna i detta parlament så är det enbart parlamentet självt som kan agera och ingen annan , för om det inte var så , så skulle europaparlamentets auktoritet och representativitet allvarligt hotas under de kommande åren och vår institution skulle inte utvecklas så som den borde .
det är minst lika viktigt att ingen skall kunna vägra lämna ut handlingar till europaparlamentet och dess utskott .
moral , disciplin och sekretess när det gäller de frågor som delegeras skall vara något som avgörs av ledamöterna i detta parlament , och inte något som bestäms utifrån av någon annan .
låt mig understryka att det inte existerar någon europeisk lag , utan ett diversifierat rättssystem i de olika medlemsstaterna .
vi löper risken att delegera frågor som rör samma brott och som sedan kommer att bestraffas olika .
jag håller med om att man bör inrätta ett undersökningssystem , men jag är lika djupt övertygad om att man måste ge rätten att försvara sig samma möjligheter och samma ställning .
jag håller inte med om att man hur enkelt som helst skall kunna göra europeiska gemenskapens tjänstemän till brottslingar : angiveri är en metod som inte hör hemma i det tredje millenniet .
avslutningsvis vill jag säga , herr talman , att från detta parlament bör utgå en tydlig signal om demokratiska principer : vi skall genomföra reformer som gör att parlamentet växer och som utvidgar dess befogenheter , inte som gör att det går tillbaka i utvecklingen .
denna debatt om van hulthens betänkande avslutar en av de mest traumatiska perioderna för de europeiska institutionerna sedan de skapades 1957 .
europaparlamentets vägran att bevilja ansvarsfrihet och den definitiva vägran att bevilja ansvarsfrihet för 1996 års budget , den misstroendeförklaring som bordlades i denna kammare av olika skäl för ett år sedan och den första rapporten från den oberoende expertkommittén om reformering av kommissionen som ledde till kommissionärernas massavgång är nu europeiska folksägner .
de av oss som var inblandade i dessa historiska händelser är väl medvetna om att inga av dessa omvälvningar skulle ha skett om vi inte hade agerat med parlamentarisk makt för att kräva förändringar i kommissionens sätt att fungera .
minns att ministerrådet , som är frånvarande igen denna debattkväll , beviljade ansvarsfrihet för 1997 - inte 1996 - samma dag som kommissionen avgick , 15 mars .
nu har vi kommit till den andra rapporten från den oberoende expertkommittén , vilken vi redan har haft tillfälle att välkomna och kort debattera i september .
det viktigaste för oss i ppe är att tillse att allmänhetens förtroende för europeiska kommissionen återställs .
ytterligare steg för att bygga ett starkt europa kommer inte att tjäna någonting till om de europeiska folken uppfattar att det inte finns något lämpligt system för demokratisk kontroll av övernitiska tjänstemän .
inte under några omständigheter kommer vi att släppa i från oss de landvinningar vi har gjort under de senaste månaderna , vilka vi tror är till gagn för öppenheten och insynen .
det bekymrar oss därför att se skurarna av tillkännagivanden från kommissionen under de senaste veckorna där kommissionär kinnock lägger olika policyförslag som skall ingå i en vitbok som snart kommer .
detta avslöjar en önskan att gå snabbt fram , men det ger också intrycket att kommissionen befinner sig i sändningsläge snarare än i lyssningsläge .
vår oro förstärks om det rykte som rapporterades för några dagar sedan stämmer - nämligen att kommissionen kraftigt vill begränsa parlamentets tillgång till information .
detta var när allt kommer omkring en av orsakerna till att den förra kommissionen föll .
har man inte lärt sig läxan ?
vetskapen om att ramen för förhållandet mellan europaparlamentet och europeiska kommissionen ännu inte är framförhandlad ledde till att vi var oense med föredraganden när vi diskuterade hans betänkande i utskottet .
vi kunde absolut inte instämma i hans åsikt att det skulle vara förnedrande för parlamentet att ta fram detaljerade instruktioner om vad vi vill att kommissionen skall ta upp i sitt reformpaket .
ju mindre exakta vi är i våra resolutioner , van hulthen , ju mer utrymme får kommissionen och era tidigare kolleger i rådet att göra vad de vill .
vi anser att det stora antalet rekommendationer i den oberoende expertgruppens rapport bör genomföras .
vi har , för ppe-de-gruppens räkning , framlagt alla rekommendationerna i expertgruppens rapport för utskottet , och många av dem har nu tagits med i betänkandet vilket helt förändrar van hulthens betänkande i utskottet .
vi har framlagt några ändringsförslag som föll i utskottet , särskilt vår önskan att uppförandereglerna skall ses över . främst vill vi lägga in hänvisningen till förtjänster och ledarförmåga som ni , herr kommissionär , när vi hade vår utfrågning i september , accepterade skulle innefattas i dessa uppförandekoder , särskilt beträffande tillsättningar och befordran .
när vi ser framåt vet vi att vi befinner oss i början av en lång process av kontinuerlig reformering av europeiska kommissionen .
vi vill särskilt se att bilden av kommissionens tjänstemän som hårt arbetande och mycket kompetenta bekräftas av yttervärlden - ett rykte som har fördunklats av ett fåtal individers olämpliga uppträdande .
herr kommissionär , ni är säkert medveten om varför krisen uppstod eftersom ni var med i den förra kommissionen .
i ett nötskal : programverksamhet bedrevs utan att det fanns tillräckliga personalresurser tillgängliga .
vi uppmanar er att ta tillfället i akt att fastställa det verkliga bemanningsbehovet för kommissionen på basis av den viktiga verksamhet den ansvarar för .
vår inställning i budgeten för 2000 var mycket klar i denna fråga .
vi kommer att vara vaksamma de närmaste fem åren för att säkerställa att de reformer som nu föreslås genomförs fullt ut och vi kommer att stödja ansträngningar att modernisera institutionerna .
men å andra sidan kommer vi inte att tveka att dra in vårt stöd vad gäller det finansiella eller annat om åtgärder skulle vidtas som inte överensstämmer med den öppenhet kommissionens ordförande romano prodi lovade innan han utsågs .
låt oss hoppas att vi kan undvika institutionella omvälvningar genom att föra en ständig dialog som från början utgår ifrån att parlamentet skall vara en jämställd partner i besluten om reformeringen av kommissionen .
herr talman ! jag måste börja med att be om ursäkt för att jag inte kan vara tillnärmelsevis så dramatisk som elles i min föredragning .
låt mig först tacka van hulthen för hans betänkande .
det skulle ha varit fel av parlamentet att okritiskt stoppa in varenda rekommendation från ett utomstående organ , för parlamentet bör ha en egen uppfattning om dessa frågor .
det är rätt att vi har ett fokuserat betänkande , vilket är vad van hulthen har producerat .
tillåt mig att uppmana elles att inte spänna vagnen framför hästen .
ja , socialisterna förlorade en hel del saker men de har inte gått igenom i plenum än och låt mig varna honom för att de kanske inte gör det i morgon .
jag skulle vilja tacka kommissionär kinnock för alla hans ansträngningar hittills .
han har varit tydlig om att han har förpliktigat sig att genomföra en radikal förändring .
försöket att skapa och införa ansvar är centralt i detta .
det är klart att detta måste utvecklas på alla nivåer och att man måste uppfatta behoven på alla nivåer inom kommissionen .
det står klart att vi behöver en förändring av budgetförordningen .
vi måste sätta stopp för att människor skyller ifrån sig på varandra .
när fel uppstår inom kommissionen måste vi ställa någon till ansvar .
vi måste få försäkringar om att konsekvent underlåtenhet att sköta sina uppgifter skall leda till avsked .
detta är naturligt på andra håll , men tycks vara ett extremt radikalt förslag när det ställs till kommissionen .
vi kan inte fortsätta med en situation där inkompetens , misskötsel och bedrägeri kostar de europeiska skattebetalarna pengar och ger dem dålig service .
jag skall ge er ett exempel på detta .
i revisionsrättens rapport för 1998 kostade en felberäkning av växelkurserna beträffande italienskt vin europas skattebetalare mellan 8 och 10 miljoner brittiska pund .
det står klart att detta inte är acceptabelt .
vad hände med den person som var ansvarig för felräkningen ?
vi behöver ett system som ger incitament och befordran och denna befordran skall ske på grundval av meriter .
vi inser att de flesta av tjänstemännen inom kommissionen arbetar extremt hårt .
men vi inser också att vissa rutiner är föråldrade .
vi ser fram emot att få läsa kommissionens hela förslag till reform och vi ser fram emot att utarbeta detaljerna jämsides med kommissionen för , trots det elles just sade , har kommissionären gjort ett åtagande att diskutera det med parlamentet före den 1 mars .
vi måste också inse att man inte skall kasta sten i glashus .
europaparlamentet har inte precis varit snövitt i sitt uppträdande under historiens gång .
vi har långt kvar innan vi är perfekta själva .
vår egen personalpolitik är förlegad .
vissa av våra arbetsrutiner behöver reformeras radikalt .
jag hoppas att europaparlamentet kommer att hålla fast vid kommissionens rockskört i denna reformprocess .
vi godkänner förslagen om verksamhetsbudgetering .
vi inser att detta innebär disciplin från kommissionens tjänstemäns sida och vi inser också att vi har ett ansvar i parlamentet för disciplin när vi talar om negativa prioriteringar .
låt mig slutligen säga att kommissionen behöver arbeta på sina relationer med allmänheten .
europas skattebetalare behöver lugnas .
kommissionens öde , hela europeiska unionens öde , beror på om denna reform kan genomföras .
detta är huvudfrågan , att dessa förslag genomförs .
herr talman ! jag skulle vilja börja med att framföra mina komplimanger till föredraganden , herr van hulten , för hans första betänkande .
jag beundrar honom särskilt för att modet inte svek honom när han drunknade i så många ändringsförslag .
jag tror att den oberoende expertkommitténs rapport har varit en nyttig rapport , och jag tror också att det är nyttigt för parlamentet - vilket också morgan sade - att vi också för en gångs skull ber expertis utifrån att se över hur vår administration sköts .
jag skulle vilja understryka ett par av de många punkterna i van hultens betänkande , det beror inte på hur pass viktiga de är utan det är helt enkelt godtyckligt .
först och främst anser jag att kommissionen måste ägna mycket större uppmärksamhet åt att bevara dokument på ett betryggande sätt .
kommissionens arkiv lämnar åtskilligt övrigt att önska .
vi lade märke till detta när vi skulle undersöka fléchard-affären som för övrigt inte på långa vägar är utredd ännu .
konstigt nog hade mycket viktiga dokument försvunnit från kanslierna , till och med från ordförandens , från olika generaldirektorat , och det är helt klart något som inte får förekomma .
om parlamentet vill göra en ordentlig kontroll måste dessa dokument vara tillgängliga , och jag skulle gärna vilja veta vad kommissionen tänker göra för att förbättra detta .
sedan något om kontrollen i efterhand , revisionsförklaringen .
det har också delvis framkommit i van hultenbetänkandet .
jag tror att det skulle vara bra om vi började ge rapportsiffror per kategori och per sektor om hur budgeten verkställs .
nu är det allmänna intrycket att allt i europa som har med budgeten att göra är dåligt .
det står klart att vi under de senaste åren sett en förbättringstendens i fråga om jordbruk och en försämrande sådan i fråga om utgifterna för strukturella åtgärder .
är det acceptabelt ?
jag skulle vilja föreslå kommissionen att fastställa en deadline för genomförandet av strukturutgifterna .
när vi antar nya medlemsstater får det inte vara så att vi ännu inte bringat ordning i eget hus .
herr talman , kolleger ! först och främst vill jag rikta ett tack till kollega van hulten .
det är hans första betänkande här i plenum .
det är värt att gratulera , även om jag naturligtvis beklagar att han inte förklarat detta betänkande på sitt eget modersmål .
bästa kolleger ! det är ett betänkande som varit svårt att få till stånd , och kanske kommer det för sent .
det har enligt min uppfattning framför allt att göra med bråket mellan de två stora grupperna i vårt budgetkontrollutskott .
låt oss vara ärliga .
den andra rapporten från den oberoende expertkommittén kom i september .
nu har det gått ytterligare fyra månader .
under tiden har van hulten drunknat i ändringsförslag , mer än 100 ändringsförslag under den första omgången .
han satte i gång på nytt , skrev om sitt betänkande , tog hänsyn till en stor mängd förslag , men möttes av ytterligare nästan 100 ändringsförslag under den andra omgången .
allt detta har således lett till , och det är jag litet orolig för , att betänkandet blivit för detaljerat , för omfångsrikt och framlagt för sent .
dessutom godkände , efter vad jag fått höra , kommissionen alldeles nyligen i dag ett förslag om reformeringen av kommissionen som kommer att skickas runt till olika institutioner för vidare konsultationer och även till vårt parlament hoppas jag .
skulle kinnock kanske vilja lyfta på förlåten redan i kväll ?
kollega van hulten ! min grupp av gröna och regionalister kommer inom kort att stödja förslagen under plenum i morgon eftermiddag om att ytterligare förbättra detta betänkande något .
det ju ingen mening med att ord för ord ta upp de många goda rekommendationerna från den oberoende expertkommittén i ert betänkande .
när vi i morgon således kommer att rösta emot vissa ändringsförslag eller emot vissa punkter är det absolut inte på grund av innehållet , utan i avsikt att göra en mer läsbar helhet av ert betänkande .
i vilket fall som helst måste det stå klart att min grupp naturligtvis fullständigt stöder rekommendationerna från den oberoende expertkommittén .
hur som helst ser jag fram emot det dokument som godkänts av kommissionen i dag .
hur som helst ser jag fram emot den vitbok som skall komma inom kort i februari .
hur som helst måste jag meddela er , herr kommissionär , att både expertkommitténs rapport och van hultens betänkande kommer att bli riktpunkter för vår grupp , riktpunkter som kommer att tydliggöra för oss om vi , ja eller nej , skall kunna hysa misstroende eller förtroende för kommissionen prodi .
som avslutning vill jag bara säga detta .
precis som i fråga om vitboken om livsmedelssäkerhet som godkändes förra veckan och släpptes till allmänheten och som innehöll en konkret tidsgräns vill vi att detta också skall gälla för den nya vitboken om reformeringen av kommissionen .
jag tror att detta är nödvändigt eftersom allmänheten ser fram emot förändring , och i vilket fall som helst vill min grupp att en tydlig förändring har förverkligats fram emot slutet av år 2002 .
herr talman ! det är bra att detta betänkande har kommit till , men det behövs egentligen mer .
bedrägeri , dålig förvaltning och svågerpolitik uppstår inte av en slump .
de får den största chansen om den demokratiska kontrollen av penningflödena är ringa .
via strukturfonderna pumpas en stor del av den europeiska budgeten runt .
det är meningsfullt endast så länge det handlar om solidaritet där rika medlemsstater bidrar till fattigare medlemsstaters inkomster och utveckling .
men det förekommer också pengar som pumpas runt och som via bryssel åter går till samma rika medlemsstater .
kommuner och regionala myndigheter ser detta som sina egna pengar , men det enda sättet för dem att få dessa pengar är genom att lägga mycket pengar och arbetsinsatser på lobbyverksamhet och förhandlingar .
efter varje oavsiktlig användning av dessa pengar , och självfallet efter bedrägeri , ljuder ropet på ännu strängare kontroll .
inte ens den allra strängaste kontroll kan lösa detta problem .
den kommer på sin höjd att leda till mer byråkrati och mindre utrymme för den lokala demokratin att vinna inflytande och mindre utrymme för medinflytande för befolkningen över val av projekt och deras innehåll .
det är bättre om dessa pengar slussas direkt från de nationella myndigheterna till de lägre myndigheterna utan att ta omvägen över europa .
vi måste någon gång under de kommande åren tänka över möjligheten att ersätta strukturfonderna med en utjämningsfond som är begränsad till budgetstöd för medlemsstater eller deras delstater med en låg inkomst per capita hos befolkningen .
det är förmodligen den enda vägen för att nå fram till mindre bedrägeri , mindre overhead-kostnader , mer öppenhet och mer demokrati .
herr talman ! det har fortfarande inte gått ett år och det är redan en uppenbar skillnad mellan det sätt på vilket parlamentet behandlar det första och det andra betänkandet .
det första betänkandet gavs omfattande publicitet , det diskuterades högtidligt och utnyttjades därefter , tillsammans med den polemik och de läckor till pressen som föregick det , till att massakrera kommissionens ordförande och därefter de flesta av kommissionärerna , trots att de inte hade något att göra med bedrägerier , tjänstefel och nepotism .
när man nu läser det som hände för knappt ett år sedan verkar det tydligt att det betänkandet skulle kunna användas till vad som helst utom att skapa klarhet eller genomföra reformer , som man hävdar i dag . på samma sätt är det sant att detta andra betänkande , som i stället skulle kunna lägga fram betydligt konkretare uppgifter , beställdes i det uttalade syftet att inte behandla specifika fall , varför det knappast är intressant att följa upp de olagligheter som nämns .
det intresserar inte de stora grupperna i detta parlament , och inte heller de flesta av de fackföreningar som i ord anstränger sig att försvara den europeiska förvaltningen , men som i själva verket bara är intresserade av att skydda sina egna medlemmar , och att därvid på ett diskutabelt vis använder de omfattande maktbefogenheter de tilldelats .
fackföreningsrepresentanter finns det i disciplinråden och i kommittén för tjänsteföreskrifterna , vilket gör det omöjligt att avlägsna de felande tjänstemännen eller att ändra på tjänsteföreskrifterna .
fackföreningsrepresentanter sitter också , obegripligt nog , i urvalskommittéerna , och jag skulle inte bli förvånad om inte företrädare för fackföreningarna också ingår i olaf , vilket gravt skulle skada denna institution som åtminstone formellt borde kunna ge garantier om att stå fri från de olika parterna .
jag förstår med andra ord varför vi träffas vid denna tidpunkt , som i regel är avsedd för annat och inte för debatt , diskussion och information .
herr talman ! när det gäller er egen reform , är kommissionen i knipa .
efter de händelser som ledde till att den tidigare kommissionen avgick , finns det en enorm förväntan .
jag får ibland intrycket att förslagen även här i kammaren får större bifall , ju mer radikala de låter .
å andra sidan kan man inte enbart med ett par penndrag ändra på förhållandena från i dag till i morgon , och svårigheterna börjar så snart det gäller genomförandet , så snart man skall tala om detaljer .
det är möjligen förklaringen till varför vi också i budgetkontrollutskottet haft fler svårigheter än väntat .
trots detta kan resultatet som det nu föreligger ses som beaktansvärt , och jag vill uttryckligen tacka kollegan van hulten för hans arbete med detta betänkande .
om detta betänkande nu inte än en gång urvattnas genom att man antar ändringsförslag , ger vi därmed kommissionen på några avgörande punkter klara och otvetydiga uppgifter .
låt mig börja med den viktigaste uppgiften .
vi vill inte avskaffa ekonomistyrningen .
det måste även i fortsättningen vara möjligt för styrekonomen att göra en granskning innan ekonomiska åtaganden eller betalningar genomförs , inte i alla enskilda fall , men alltid där det finns osäkerhet eller risker .
här ger kommissionen fel signaler , till exempel när man döper om generaldirektoratet för ekonomistyrning till generaldirektorat för revision .
kommissionens organisationsschema går väl lätt att ändra , men det blir svårare när kommissionen angriper lagtexterna , i synnerhet budgetförordningen .
jag har inte räknat efter så noga , men gemenskapens budgetförordning och de dithörande genomförandebestämmelserna talar på nästan 100 olika ställen om styrekonomen , hans oberoende och de uppgifter han har .
detta kan inte ignoreras eller kringgås , inte heller med s.k. soft law , som det en gång antyddes under ett sammanträde med vårt utskott .
oberoende av sådana rättsliga överväganden vore det också med tanke på sakens natur ett oförlåtligt fel att avskaffa ekonomistyrningen i dess klassiska bemärkelse just i det ögonblick , när de i kommissionen som är ansvariga för detta äntligen inte längre står helt ensamma , utan kan bli ett led i en kedja av fungerande kontroll- och undersökningsmekanismer .
vår idé är att det i framtiden skall vara tre mekanismer som griper in i varandra , den oberoende förhandskontrollen som görs av styrekonomen , den åtföljande efterhandskontrollen som görs av den interna granskningsenhet som skall inrättas , även kallad revisionstjänsten , och slutligen det målinriktade uppspårandet av oriktigheter som görs av olaf , den nya byrån för bedrägeribekämpning .
det är bra att kollegan van hultens betänkande framställer sammanhanget mellan alla tre områdena och också klargör var de avgörande brister ligger , som skall åtgärdas .
helt kortfattat vill jag säga : de disciplinära förfarandena fungerar inte , i synnerhet när det gäller att hålla tjänstemän till räkenskap för sitt olämpliga uppträdande även ekonomiskt .
det finns en stor gråzon och många oklarheter i fråga om de straffrättsliga påföljderna , och just här är det som vi har hört från kommissionen , snarast vagt .
jag kan bara understryka att detta är de verkligen hårda nötter som äntligen måste knäckas !
herr talman ! först och främst vill jag helhjärtat gratulera min kollega van hulten .
det är roligt att kunna säga att han kommer från vår delegation , och jag tror att jag kan få vara litet stolt över honom .
hur som helst vill jag gratulera honom till hans betänkande .
herr talman ! kommissionens avgång har också skapat en kultur som kännetecknas av rädsla hos många tjänstemän i hierarkin och den stora byråkratin .
hela pläderingen om att förändra kulturen till en ansvarskultur förefaller mig vara mycket grundläggande .
jag har i utskottet utveckling och samarbete på mycket nära håll kunnat uppleva hur tusentals projekt stagnerat , att ibland 80 procent av pengarna inte kommer till användning , att ibland en enorm damm av pengar uppstår , inte på grund av det faktum att pengarna inte är helt nödvändiga , inte på grund av det faktum att det inte finns några goda förslag , utan på grund av att hela systemet i sig självt har låst sig .
brist på ansvar , alldeles för mycket ex ante , alldeles för lite ex post och därför alldeles för litet kultur som kännetecknas av verkligt effektiv förvaltning .
det vore fantastiskt om vi med detta betänkande skulle kunna ge signalen till resultatinriktad förvaltning och organisera hela arbetet på grundval av denna .
jag hoppas verkligen på att den insats som vi har gjort här , när kommissionens preliminära rapport blir den officiella rapporten inom kort den 1 mars , kommer att bidra till att vi här verkligen kommer att få se denna förändring .
det skulle verkligen vara att göra den europeiska allmänheten en tjänst , herr talman , utan någon som helst tvekan , och genom de resultat som vi visar skulle vi också återvinna och återförvärva något av det som vi under de gångna åren uppenbarligen har förlorat .
det är det bästa stöd vi kan ge den europeiska demokratin .
om vi därmed kommer bort ifrån 50-talskulturen och övergår till nästa århundrade , då får vi här uppleva ett mycket vackert ögonblick .
herr talman ! först skulle jag vilja framföra gratulationer till michiel van hulten för hans första betänkande .
det var en tuff nollning , men i nederländerna har vi ett passande talesätt : &quot; det snabbaste sättet att lära sig simma är att direkt kasta sig ut på djupt vatten . &quot; ärade kollega !
jag tror att ni efter denna prövning skulle kunna kvalificera er till olympiska spelen .
det finns två punkter som enligt min och eldr : s uppfattning förtjänar särskild uppmärksamhet .
för det första gäller det kommissionärernas individuella ansvar .
detta måste regleras under regeringskonferensen .
vi vill dock inte att denna viktiga fråga skall komma att ligga helt och hållet i rådets händer , och därför har vi lagt fram ett ändringsförslag där vi ställer frågan om inte ett interinstitutionellt avtal skulle kunna komma till stånd mellan kommissionen och parlamentet för att sörja för att vi har en sorts fall back-position och inte lägger vår lott helt och hållet i rådets händer .
den andra punkten , vilket också min kollega mulder sagt , är att eldr anser att även europaparlamentet måste synas av oberoende experter .
detta kommer att ge ett mycket stort bidrag till att återställa de europeiska medborgarnas förtroende för denna institution .
vi kan inte vara någon trovärdig motpart till denna kommission så länge vi inte också rannsakar våra egna samveten och bringar ordning på torpet även i europaparlamentet .
det är bara om alla europeiska institutioner reformeras som vi kan få det öppna , demokratiska och handlingskraftiga europa som våra medborgare nu äntligen förtjänar .
herr talman ! även jag vill gratulera min kollega van hulten till det första betänkande han lägger fram här i parlamentet .
jag är säker på att han kommer att ha nytta av detta , bland annat i form av ett andra ännu smidigare betänkande och i en allt starkare strävan efter alla gruppers samtycke .
vid det här laget får den process med en reform av kommissionen som krävs av medborgarna inte skjutas upp längre .
i det här parlamentet har vi vid flera tillfällen , även av kommissionens ordföranden , fått ta del av deras önskan om en reform .
nu verkar det som att det skall bli allvar .
sedan en kommission har avgått och en expertkommitté har påvisat ett oräkneligt antal brister , verkar det löfte som prodi avlade den 14 september rimligt om att han inför parlamentet skall lägga fram ett fullständigt reformförslag i februari månad .
parlamentet ser fram emot ett sådant fullständigt reformprogram .
syftet med det betänkande som vi diskuterar i dag är att ge politiskt stöd till en stor del av rekommendationerna från den expertkommitté som parlamentet anlitat .
prodi har sagt att han hur som helst kommer att agera , att han föredrar att lyckas , men att rädslan för att misslyckas inte kommer att hindra honom från att agera .
därför kräver vi ett djärvt program , och i sådant fall garanterar jag att parlamentet kommer att stödja kommissionen i denna reformprocess .
vi vill ha en stark kommission som kan uträtta sitt arbete på ett oberoende och neutralt sätt , men med politiskt omdöme .
kommissionärerna bör inte betrakta sig själva som höga tjänstemän utan som verksamma politiker .
betänkandet medger deras rätt att vara aktiva politiker och tillhöra politiska grupperingar inom ramen för sitt parti .
kanske är inte det som rör befattningarna helt i sin ordning .
jag känner inte helt till er bedömning i det fallet , herr kinnock , men det är självklart att vi vill ha kommissionärer som är politiskt starka med ett politiskt engagemang .
och vi vill ha en struktur som medger en effektiv användning av varje euro , för vid varje bokslut framgår att så inte är fallet .
av den anledningen , herr kommissionär , uppmuntrar vi prodi att komma hit med ett djärvt program , och han kommer att upptäcka att han får problem med sådana grupper som riskerar sin status quo , däremot inte med parlamentet som förväntar sig djupgående och djärva förändringar .
herr talman ! jag vill tacka van hulthen för hans betänkande och säga att jag röstade för det .
så jag tar upp de saker jag inte är överens om .
jag instämmer inte i avsnitten som gäller parlamentet .
detta betänkande handlar om kommissionen .
parlamentet är ett annat ämne .
det finns ingen anledning att dra in parlamentet i diskussionen om kommissionen .
dessutom är det frågan om tax-free .
detta användes emot kommissionen av de tax-free-lobbyister som var emot det faktum att kommissionen avskaffade tax-free-försäljningen på flygplatser .
den är inte heller värd att tas in i detta betänkande .
största delen av betänkandet handlar om ekonomisk kontroll .
detta är rimligt eftersom det kommer från budgetkontrollutskottet .
men vi bör inte ge intryck av att stora summor av de europeiska resurserna sätts på spel till följd av vårdslöshet i europeiska kommissionen .
trots allt är det bara 1 procent av bnp jämfört med nationella utgifter .
vi har gått igenom allt detta förr , men en del i detta parlament är unga och verkar inte förstå hur små europeiska unionens ekonomiska medel är och att medlemsstaterna gör av med 80 procent av dessa medel .
så vårdslöshet med hur pengar spenderas inom kommissionen riskerar inga stora penningsummor .
vi måste få perspektiv på detta .
detta är någonting som man måste komma ihåg .
europeiska kommissionens verksamhet handlar till väldigt liten del om att göra av med pengar .
de har väldigt litet av den varan .
de har ett mycket större ansvar .
detta större ansvar gäller att sköta miljö , livsmedelssäkerhet , utrikeshandel , den inre marknaden och så många andra ansvarsområden som vi har gett dem utan resurserna att ta itu med dem .
jag tillhör inte dem som håller med om att det finns en stor brist på förtroende .
om det gör det är det vi i detta hus som har skapat den under det senaste året .
jag har varit här i 20 år och upplevt ett absolut förtroende mellan rådet , kommissionen och parlamentet .
vi har haft våra problem och erkänt svårigheter , men det har inte funnits något läge då medborgarna i europeiska unionen har misstrott , tvivlat på och fruktat denna byråkratiska kommission för att den har misskött våra affärer .
detta är en enorm överdrift av vilka svårigheterna var .
denna kommission borde inte för alltid behöva leva i skuggan av de misstag som ledde till att dess företrädare avgick .
även om det förekom problem - som vi måste lösa mot bakgrund av utvidgningen till exempel - överdriver vi ibland det negativa .
herr talman ! låt mig tacka föredraganden för hans utmärkta betänkande .
jag hoppas att kommissionen kommer att använda det under sitt reformarbete .
reformprocessen har nu pågått en tid och det verkar råda ett slags undantagstillstånd i kommissionen .
förvaltningen inom kommissionen fungerar helt enkelt inte särskilt bra .
det finns naturligtvis bra och duktiga anställda vid kommissionen , de flesta är det .
men vi behöver en genomgripande reformering .
det är för litet handling och för mycket onödig byråkrati .
folk skall ha tydliga befogenheter att fatta beslut , och så skall de också ansvara för dem .
budgetförordningen skall ändras .
vi är överens om att vi skall utöva en bättre kontroll av pengarna .
kommissionen och expertkommittén vill helt avskaffa förhandskontrollen .
det måste vi se upp med .
vi måste behålla en viss form av förhandskontroll av pengarna .
det räcker inte med att bara tillämpa stickprovskontroll , när pengarna betalts ut .
då kan för många oegentliga projekt smita igenom .
vi måste i stället reformera och decentralisera kontrollen .
kommissionen har inte tillräckligt med personal .
vi måste i egenskap av parlamentariker ha mod att förklara för våra regeringar och väljare i våra hemländer , att personalresurserna helt enkelt inte är tillräckliga för de uppgifter som kommissionen har att utföra .
och kommissionen skall ha möjlighet att säga nej till nya uppgifter om den inte får mer personal .
personalsystemet är för stelt .
det måste vara en större rotation av anställda , särskilt i toppen av hierarkin .
det måste också vara mycket enklare att avskeda odugliga och inkompetenta anställda .
jag är därför mycket glad över att det sker en reformering av det disciplinära förfarandet .
de mycket dåliga erfarenheterna rörande de disciplinära fallen visar ju allt för tydligt hur viktigt det är att vi genomför en reformering .
herr talman , värderade kommissionärer ! först kan jag inte låta bli att reflektera över att detta är en i stort sett nederländsk-brittisk-skandinavisk debatt vad gäller talarna .
kanske är detta litet oroande .
jag hoppas , som så många andra , att undantagstillståndet i relationerna mellan kommissionen och parlamentet är på väg bort .
vi måste komma ifrån att vi rusar iväg och släcker en brand i ett hörn för att sedan rusa vidare för att släcka nästa .
vi måste i stället , som blak sade , bygga upp ett system med klara roller .
för det första behöver vi ett hårt regelverk , som kan tillämpas .
det räcker inte med uppförandekoder och etiska kommittéer .
det måste finnas hårda regler som bland annat anger vad som kan decentraliseras , vad som kan läggas ut och vad som är oberoende .
jag tycker att det är litet oroande att man i denna debatt ropar på oberoende utan att definiera oberoende i förhållande till vad och med vilken beslutsrätt .
vi behöver alltså ett grundläggande administrativt regelverk för eu , för dess institutioner och för eu i dess relationer till medlemsstaterna .
detta saknas .
vi har efterfrågat en åklagarmyndighet och en straffrätt , men vi behöver också en förvaltningsrätt för eu .
vi skulle komma en bra bit på vägen om kommissionen antog ombudsmannens förslag till uppförandekod för god förvaltningssed som ett bindande regelverk .
van hultenbetänkandet är ett steg i rätt riktning , men det är inte tillräckligt .
för det andra måste vi också klarlägga våra egna revisionsroller .
revisionsrätten skall göra en kontroll av huruvida någonting är oförenligt med regelverket , men den skall inte kontrollera ändamålsenligheten .
det är europaparlamentet som gör den politiska utvärderingen .
vi jagar inte bovar - det får olaf göra .
säg mig vilket nationellt parlament som exempelvis får alla förundersökningshandlingar !
med den drucknes envishet vill jag också säga att offentlighetsförordningen måste bli klart bättre än de utkast som har cirkulerat på internet , annars kommer vi ingen vart i den kampen .
herr talman ! jag skulle vilja framföra ett hjärtligt tack till föredraganden för hans betänkande .
jag är glad att jag nu kan tilltala honom på nederländska , nu när även van den berg gjort detta .
annars hade jag kanske känt mig lite skyldig för det .
jag skulle vilja säga att detta betänkande har genomgått en mycket stor förbättring , även genom ändringsförslagen .
jag kommer från utskottet för sysselsättning och socialfrågor , och en föredragande hos oss är alltid stolt över att få 100 ändringsförslag , för då vet han att det är ett intressant ämne som han har tagit upp .
jag tror att det är fallet här också , men enligt min uppfattning är det en smula överdrivet att prata för mycket om dessa 100 ändringsförslag .
jag vill vidare peka på att vår samordnare i budgetkontrollutskottet är pomés ruiz som är spanjor och som således har gett ett mycket viktigt spanskt bidrag till denna debatt .
herr talman ! jag anser att en av viktigaste sakerna som nämnts är föredragandens förslag om en oberoende permanent kommitté för normer för det offentliga livet .
ett mycket viktigt förslag .
men jag är mycket förvånad över att den socialistiska gruppen vill skjuta ihjäl det förslaget genom ett förslag av morgan , för hon vill avlägsna det helt och hållet .
jag förstår inte alls hur det kan vara möjligt .
vi får å ena sidan allehanda lovyttringar ämnade för föredraganden , men samtidigt vill morgan på den här punkten , liksom på andra viktiga punkter för övrigt , litet grand följa den brända jordens taktik , vilket egentligen leder till att innehållet i detta betänkande helt och hållet försvinner .
jag vet inte om det är för att tillmötesgå kinnock . men jag känner kinnock .
kinnock vill gärna höra vad vi vill och är också fullt beredd att förirra sig bort från detta om han anser det nödvändigt .
jag anser att en sådan långtgående brända jordens taktik egentligen inte behövs .
slutligen , frågan om tjänstemännen .
jag är egentligen inte alls överens med haarder .
jag är överens om att akten om tjänstemännen egentligen har fått ett innehåll som är helt otillräckligt .
för det första läggs ingen tonvikt vid vikten av en offentlig förvaltning i största allmänhet .
för det andra nämns allehanda förslag där man måste ställa sig frågan om de nu är så förståndiga och om de kommer ge anledning till förbättring .
till exempel , vi sysslar med dessa kontor för tekniskt bistånd , och det är en viktig punkt , och samtidigt vill vi avskaffa kommissionens tillfälliga personal .
detta ligger på kollisionskurs , och jag förstår verkligen inte hur ett sådant förslag har kunnat läggas fram .
herr talman ! sedan platons republik har västvärlden systematiskt försökt ersätta folkregeringar med expertregeringar .
vårt parlament inbjöd först experterna för att hjälpa till att utvärdera europeiska kommissionens arbete och dessa utnyttjade inbjudan för att ta dess öde i sina händer .
i denna andra rapport har experterna redan tagit ett nytt steg och kritiserar de politiska grupper som i parlamentet tvekade att avsätta europeiska kommissionen , på grund av det gemensamma politiska medlemskapet med några av dess medlemmar , och anser att detta problem övervinns genom att förbjuda kommissionärerna att tillhöra politiska grupper .
enligt experterna borde parlamentet inte ha kontrollmakten över europeiska kommissionen och borde i denna uppgift ersättas av en permanent och inte vald kommitté för normer för det offentliga livet , vilken förmodligen skulle bestå av en annan grupp experter .
i denna andra rapport lär experterna oss att italien finansieras av sammanhållningsfonden , att europeiska regionala utvecklingsfonden och socialfonden utgör två tredjedelar av strukturfonderna , att additionalitets- och komplementaritetsprinciperna i strukturfonderna är likvärdiga , att jordbrukslobbyn ålägger garantisektionen inom europeiska utvecklings- och garantifonden för jordbruket ( eugfj ) finansieringen av landsbygdens utveckling , och att samarbetsprincipen bara tillämpas på kommissionen och medlemsstaterna .
denna visdom är 100 procent ideologi och 0 procent kunskap .
det är inte på det sättet vi stöder reformen av de europeiska institutionerna med full respekt för de demokratiska institutionerna .
hultenbetänkandet var inledningsvis ett lysande betänkande och jag vill ge min djupa och innerliga hyllning till det som har gjorts här av vår kollega hulten .
tyvärr förändrades det undan för undan i sämsta möjliga riktning , och gjordes om till ett dokument som faktiskt försvarar något vi inte kan acceptera .
herr talman , herr van hulten ! ert betänkande har gjort sig förtjänt av följande adjektiv : vågat , krävande , komplext och jag tror att det är viktigt för ett första betänkande .
ta därför det jag nu kommer att säga som kritik för motsägelsens egen skull , något jag tror kan vara berikande för denna debatt .
jag uppfattar detta betänkande som onödigt ordrikt , långrandigt , rörigt och oklart vad beträffar de idéer som framförs .
onödigt ordrikt kanske är det värsta adjektivet , och ni är inte ansvarig för detta , utan det ansvaret åligger parlamentet .
det vill säga , om parlamentet ger i uppdrag åt en expertkommitté - och jag skall inte upprepa det casaca sade , men jag håller med honom - att analysera ett problem , vad är det då för mening med att ge sig in på en medeltida tradition som innebär att tolka uttolkarna och så vidare ad infinitum .
det är uppenbart att vi väntar på en reform av kommissionen , vi väntar på de förslag som kommissionen kommer att lägga fram , och parlamentet bör sedan uttala sig om dessa .
bland annat måste vi ge uttryck för vårt förtroende för kommissionen .
långrandigt .
jag skall inte nämna hur pass omfattande detta betänkande är .
jag vet inte om det slår rekord bland alla de resolutioner som har framförts här , men det gör det åtminstone bland denna typ av resolutioner .
jag tror inte att vi tidigare har haft någon resolution - och då bör man tänka på att vi ger upphov till omfattande resolutioner här i parlamentet - som har innehållit stycken med mer än 16 rader utan punkt .
dessutom är det rörigt .
jag skall inte upprepa det man redan har sagt beträffande analysen av frågor som rör parlamentet .
denna borde bli föremål för ett annat betänkande och det måste vi se till , och det är viktigt att vi funderar över detta , men inte inom ramen för detta betänkande .
och slutligen , herr talman , skall jag inte gå in på några exempel , men ärligt talat förekommer det flera sådana där det juridiska språket används med en oroväckande brist på exakthet .
därför - så här sammanfattningsvis - ser jag fram emot - vi är många som ser fram emot -er rapport , herr kommissionär kinnock , så att vi kan uttala oss för denna , vilket är det som parlamentet bör göra .
herr talman ! av omfånget och detaljflödet i förslagen till nödvändiga reformer kan man sluta sig till vikten av en sådan reform .
men med tanke på de händelser som har utlöst dessa ansträngningar , är nödvändigheten också uppenbar .
förhoppningarna och förväntningarna har blivit så mycket större på grund av de starka tillkännagivandena av kommissionärerna prodi och kinnock i kammaren och i budgetkontrollutskottet .
i betänkandet lägger man särskilt märke till begreppet öppenhet .
att garantera denna är en huvudfråga .
vikten av fullständigt föreståeligt arbete kan heller inte påpekas ofta nog .
men det handlar inte enbart om en byråkratisk reform , utan snarare om att demonstrera den goda viljan gentemot våra medborgare .
deras förtroende för eu : s politik måste vinnas tillbaka .
medborgaren begär snabb och öppen tillgång till institutionen och till läsbara föreskrifter .
hans förståelse beror av detta , och han vill ha en framgångsrik politik och uppfattar detta samtidigt som en självklar tjänst åt den myndiga medborgaren .
om reformen skall lyckas beror till väsentlig del på kommissionens egna initiativ .
men det irriterar mig när jag i dag hör att kommissionen nu säger att den bara vill diskutera delrapporten informellt med parlamentet .
men ert föredrag , herr kinnock , i budgetkontrollutskottet kommande tisdag får inte bara vara enkelriktat , utan vi som parlamentariker vill och måste vara med om utformningen . och det ligger också utanför min politiska förståelse när det denna vecka äger rum ytterligare en presskonferens innan vi i det ansvariga budgetkontrollutskottet noggrant har diskuterat förslaget .
jag tror , herr kinnock , trots all personlig framgång , att kommissionen måste göra en hel del mer för att uppfylla våra berättigade höga förväntningar .
fredsprocessen i mellanöstern ( fortsättning )
nästa punkt på föredragningslistan är fortsättningen på debatten om rådets och kommissionens uttalande om fredsprocessen i mellanöstern .
) herr talman ! vi förstår kommissionär patten mycket väl .
jag vill bara säga att förbindelserna med madrid i vanliga fall är ganska så bra , och att jag därför snart hoppas få se honom där .
de uttalanden vi under dagens lopp har hört om fredsprocessen i mellanöstern kommer mycket lägligt efter den pressande rundresa minister gama - jag beklagar hans frånvaro - tillsammans med tre andra representanter från rådet gjorde i området .
de nyheter man rapporterat om i massmedia skulle kunna få oss att se pessimistiskt på situationen .
jag tror ärligt talat att en utvärdering av det här slaget inte överensstämmer med verkligheten .
jag delar därför kommissionär pattens positiva inställning .
jag skall förklara varför : det är sant att den israeliska regeringen har flyttat fram det tredje överlämnandet till de palestinska myndigheterna av mark på västbanken .
men det är också sant att man sedan sharm el-sheikh har överlämnat 39 procent av västbanken och två tredjedelar av gazaremsan till palestina och att - vilket är än viktigare - nämnda avtal fram till nu har följts till punkt och pricka , till och med uppskovet är ett prerogativ från den israeliska regeringens sida som förutsetts i sharm el-sheikh .
förutsatt , givetvis , att det inte dröjer mer än tre veckor , vilket är vad premiärminister barak har lovat .
å andra sidan är beslutet att flytta fram den andra samtalsrundan , som inleddes i shepherdstown av arabrepubliken syrien , tvivelsutan en viktig händelse , men jag är övertygad om att hoppet från den 3 januari inte kommer att gå förlorat .
herr talman , det faktum att kammarens alla politiska grupper inställer sig till den här debatten , som alltid är kontroversiell , med ett resolutionsförslag som man enhälligt har bifallit tycker jag är avgörande för vår politiska vilja att bestämt stödja de pågående fredsförhandlingarna .
med samma kraft tar vi avstånd från våldshandlingar för att lösa meningsskiljaktigheter , må vara djupa , parterna emellan .
enligt min mening är detta en garanti för båda parter , såväl ur politisk som ekonomisk synpunkt , för de åtaganden som kan förväntas av europeiska unionen när det gäller kostnaderna för den fred vi alla så hett eftertraktar .
för att kunna garantera säkerheten i området och för att kunna bidra till att mildra rådande sociala skillnader förnekar ingen att detta är absolut nödvändigt .
men det uppmärksammar också europeiska unionens krav på att politiskt få delta i processen , i enlighet med vårt ekonomiska stöd så att det offentliggörs på motsvarande sätt , eftersom inte heller vi gör anspråk på att vara bankirer .
europaparlamentets ordförande och hennes kommande resa till området kommer tvivelsutan att bidra till detta .
herr talman ! jag vill tacka kommissionär patten för en utförlig beskrivning .
jag vill gärna säga att jag ansluter mig till den ton som galeote quecedo angav här .
vi i parlamentet stöder starkt fredsprocessen i mellanöstern .
det är ju en fredsprocess som äntligen är på gång .
trots svårigheter och förseningar , är det ändå en skillnad som mellan natt och dag om vi tänker på hur processen såg ut för ett år sedan .
för det första innehåller sharm el-sheikh-avtalet en konkret tidsplan som alla vet för genomförandet av israels åtaganden ; det gäller då interimsavtalet samt hebron- och wye-avtalen .
medan förhandlingarna om slutlig fredsuppgörelse har inletts , tror jag att det är viktigt att hålla isär de två .
brist på framsteg i slutstatusförhandlingarna bör inte äventyra genomförandet av de tre ovannämnda interimsavtalen .
vad vi behöver bevaka i detta sammanhang är hur det går med hamnen i gaza , den nordliga transitrutten mellan gaza och västbanken , ytterligare frisläppande av säkerhetsfångar och genomföranden av de ekonomiska åtagandena .
den andra punkten gäller syrien .
där är naturligtvis gränsfrågan central .
hur förhandlingarna går där , vet vi inte ännu .
det viktiga är emellertid att de har inletts .
en viktig fråga i sammanhanget är den framtida vattenfördelningen .
golan svarar i nuläget för mellan en tredjedel och en sjättedel av israels vattenförsörjning .
den tredje aspekten är fredssamtalen i syrien som är nära sammankopplade med frågan om israeliskt tillbakadragande från södra libanon .
enligt uppgift från unifil , finns det nu konkreta tecken på att israel förbereder ett tillbakadragande , vilket vi välkomnar .
utestående tvistefrågor är naturligtvis även där vattenproblematiken och de libanesiska palestinaflyktingarnas situation .
min sista punkt gäller den kommande palestinska staten .
den kan komma att utropas under detta år , med eller utan israels stöd .
regeringen barak har låtit förstå att man är inställd på att sluta ett fredsavtal med en stat som motpart .
även om inte förhandlingarna är avslutade i september detta år , finns det inga fördragsmässiga hinder mot att en palestinsk stat skall utropas efter detta datum .
i detta sammanhang är det då viktigt för oss som stöder tanken på detta , att det blir som kommissionär patten sade , nämligen en stat med insyn och att det blir en demokratisk stat .
det vill vi alla medverka till .
jag skulle gärna först och främst vilja hänvisa till den gemensamma resolution som skall läggas fram som avslutning på den här debatten och till vilken min grupp bidragit och som vi naturligtvis godkänner .
mer specifikt vill jag dock uttrycka min glädje över att israel och syrien efter så lång tid återigen samtalar för att lösa sina meningsskiljaktigheter .
de nya förhandlingarna är i alla fall ett viktigt steg mot en varaktig fred i mellanöstern .
därför är det synd att de här fredssamtalen skjutits upp tills vidare .
båda parter kommer mycket riktigt att behöva göra stora insatser .
en varaktig fred i det här området kan förverkligas först genom ett avtal i vilket säkerheten för de israeliska gränserna och syriens integritet kan garanteras .
för det behövs också fasta diplomatiska förbindelser och en oavbruten dialog .
förutom de bilaterala mötena med syrien hoppas jag att israel inom överskådlig tid även skall inleda förhandlingar med libanon och att en multilateral process skall visa sig möjlig inom ramen för det ekonomiska och regionala samarbetet .
det är ändå beklagansvärt att europeiska unionen , en av de viktigaste ekonomiska givarna , fortfarande inte kan spela en viktig politisk roll i fredsprocessen .
den här fredsprocessen i mellanöstern är en av prioriteterna för europeiska unionens gemensamma utrikes- och säkerhetspolitik .
här har solana , den höga representanten i rådet , en särskild funktion .
kommissionen och medlemsstaterna måste också uppmuntras att stödja projekt som kan hjälpa till att bygga upp förståelse och partnership mellan de olika folkgrupperna i det här området .
jag måste också påpeka barcelonaprocessens betydelse som ju måste ha ett positivt inflytande på det regionala samarbetet .
i det avseendet stöder vi libyens deltagande , på villkor att landet erkänner de mänskliga rättigheterna , avstår från att ge stöd till terrorister och ger sitt fullständiga stöd till fredsprocessen .
det kvarstår naturligtvis många olösta problem och obesvarade frågor , även med palestinierna .
alla vet att fredsprocessen är en lång och tung process men vi är övertygade om att med nödvändig tillförsikt , med den oumbärliga politiska viljan och med den ihärdighet som behövs så kommer vi att nå vårt gemensamma mål , nämligen ett fredligt och välmående mellanöstern .
herr talman ! det är glädjande att fredsförhandlingarna , trots vissa uppskov och problem , pågår såväl mellan israel och palestina som mellan israel och syrien .
sanningens minut närmar sig .
är israel berett att följa fn : s resolutioner och återlämna de arabiska områden som erövrades 1967 i utbyte mot fred och säkerhet ?
kommer israel att låta palestinska flyktingar återvända eller få kompensation ?
kommer israel att dela med sig av jerusalem och floden jordans vatten ?
kommer det fria palestina att bli en fullt demokratisk stat och därmed pålitlig som fredspartner ?
kommer syrien att fullt ut acceptera israels existens och införa demokrati och rättsstatlighet ?
att huvudansvaret för fredsprocessen ligger på ockupanten israel hindrar inte att också de arabiska parterna har ett stort medansvar .
mellanösternfreden angår oss emellertid alla .
därför är det bra att eu agerar som fadder till den palestinska staten .
mot denna bakgrund vill jag avsluta med en märklig historia i eu-landet sverige . där hålls en internationell regeringskonferens om hitlers judeutrotning , vilket självklart är ett välkommet initiativ .
bland fyrtiosju inbjudna stater från samtliga världsdelar finns emellertid inte en enda av de arabstater som ingår i eu : s barcelonaprocess .
detta har tolkats som att den arabiska hållningen gentemot israel av européer skulle betraktas på samma sätt som nazismens antisemitism , vilket ju är fullständigt felaktigt .
arabvärldens israelkritik har byggt på samma sorts antikolonialism som exempelvis algeriets frihetskamp mot frankrike .
men i dag har ju egypten , jordanien och palestina fördragsfäst fred med israel .
därför undrar jag om inte kommissionär patten håller med mig om att det hade varit rimligt och lämpligt att åtminstone någon arabstat hade varit inbjuden till förintelsekonferensen i stockholm .
herr talman ! jag vill verkligen tacka kommissionär patten för de kunskaper han gett prov på när det gäller svårigheterna i fredsprocessen och den utmaning som europeiska unionen har antagit när det gäller att förverkliga den .
det är verkligen dags för fred i mellanöstern .
det är dags att avsluta den epok i historien som inleddes med balford-förklaringen 1917 och det arabisk-israeliska kriget 1948 .
det är dags att det äntligen blir säkra gränser för samtliga länder i området , politiska , sociala och ekonomiska rättigheter , mänskliga rättigheter som erkänns och tillämpas i syrien , palestina och israel , överallt .
det handlar också om att varje folk och varje individ skall kunna leva självständigt och demokratiskt , men för att det skall kunna förverkligas är det nödvändigt att samtliga parter i konflikten har modet att tillämpa fred och rätt , att man erkänner den andre som en partner och inte som en undersåte som man måste bevilja eftergifter .
jag tänker i första hand på knuten palestina-israel , men det gäller även de områden som ockuperades i golan 1967 och den södra delen av libanon efter 1982 .
israel måste ta sitt ansvar , lämna de ockuperade områdena och dela på vattenresurserna , men samtidigt måste israel få garantier för sin säkerhet och kunna leva i fred i ekonomiskt och politiskt utbyte med samtliga länder i området .
men säkerheten gäller inte bara israel .
samma sak gäller de övriga länderna , i första hand palestinierna som fortfarande lever under militär ockupation och som fortfarande i dag , trots de avtal som undertecknats från och med oslo , ser sin mark konfiskerad i områdena b och c. efter oslo och fram till och med den 17 oktober 1999 har 174 tusen dunans mark konfiskerats , varav 8 462 under den nya regeringen barak .
träd har ryckts upp med rötterna , hus har förstörts och framför allt i östra jerusalem har utnyttjandet av vattnet inskränkts eller förvägrats , medan bosättningarna fortsätter och hela tiden ökar .
det råder emellertid inget tvivel om att i och med att den nya regeringen valts så har framsteg gjorts , åtminstone har man börjat förhandla igen .
men det kan inte finnas någon stabil och varaktig fred i mellanöstern om inte palestinierna får sin egen stat , om de inte fritt kan röra sig på sitt eget territorium .
det internationella samfundet måste helt enkelt tillämpa resolutionerna nr 332 , 248 , 245 och 194 .
det är oroande att förbindelserna med syrien har skjutits på framtiden , liksom baraks beslut att skjuta upp tillbakadragandet av den israeliska armén och avtalen från sharm el-sheikh .
det är utomordentligt viktigt att europeiska unionen kan spela en politisk roll i förhandlingarna parallellt med sin roll när det gäller ekonomiskt bistånd .
vi kan inte nöja oss med att stå i kulisserna , vi måste i stället spela en huvudroll , utan att för den skull hamna på kollisionskurs med usa , som minister gama påpekade .
herr talman ! låt mig först uttrycka mina tack och min uppskattning till kommissionär patten för hans kommentarer här i dag , särskilt i samband med europeiska unionens roll i fredsprocessen och för att han bekräftar att vår roll inte bara innebär att vara &quot; bank &quot; för hela verksamheten .
jag blev djupt besviken när jag fick höra nyheterna i veckan om att fredssamtalen mellan israel och syrien hade skjutits upp .
jag hoppas verkligen att man kan nå en kompromiss , så att fredssamtalen snabbt kan återupptas .
vi kan emellertid inte förneka att det skett en del positiva politiska framsteg i mellanöstern under den senaste tiden .
det faktum att den syriske utrikesministern och den israeliske premiärministern nyligen satt vid samma bord i förenta staterna för första gången någonsin är ett tecken på går att övervinna det gamla hatet och fientligheterna .
de politiska ledarna måste visa verkligt mod för att anta en gemensam ram som kan leda fram till en övergripande fred i mellanöstern .
jag vet att om det går att nå ett avtal mellan syrien och israel , kommer israels premiärminister att möta verkliga protester mot alla nya avtal med syrien i framtida folkomröstningar .
bosättarna på golanhöjderna kommer att kräva kompensation och det måste bli garantier rörande säkerheten .
om syrien skulle vara redo att ta itu med säkerhetsfrågan , skulle utsikterna för en lösning på israel-syrienfrågan vara goda .
vad gäller palestinafrågan inser jag att det fortfarande finns vissa svårigheter rörande genomförandet av vissa aspekter av wye-avtalet .
de största problemområdena omfattar för tillfället omstrukturering , såväl som överflyttning av territorier .
den låga graden av frisläppande av palestinska fångar och det faktum att den israeliska regeringen verkar stoppa tillämpningen av byggnadstillstånd som redan beviljats , såväl som att inte utfärda nya , utgör ytterligare hinder .
dessa frågor har uppenbarligen hejdat framstegen i förhandlingarna om den permanenta statusen , även om - tror jag - dessa samtal inte kommer att stoppas för evigt .
den största svårigheten just nu när det gäller att få igång förhandlingarna , verkar vara att palestinierna vill att man först och främst skall lösa gränsfrågan , medan den israeliska regeringen säger att denna endast kan lösas om man först når en lösning i frågan om bosättningarna och säkerheten .
för tillfället verkar det som om båda sidor har accepterat att man inte kan komma överens om någonting , förrän man kommit överens om allt .
medan , sammanfattningsvis , andra länder i mellanöstern haft betänkligheter rörande fredsprocessens allmänna riktning , nu när den syriska regeringen också deltar i fredsprocessen , är egypten och andra länder i regionen redo att gå vidare .
jag hoppas verkligen att - när det gäller att förbättra säkerheten och livskvaliteten för folken i mellanöstern - alla tongivande parter så snart som möjligt ser till att ingå ett övergripande avtal om alla viktiga frågor som behöver få en lösning .
herr talman , ärade kolleger ! de olika resolutionsförslag som lagts fram i parlamentet ger en god bild av läget i mellanöstern .
det finns de som applåderar nya avtal mellan israel och syrien , men bara någon enstaka riktar uppmärksamheten mot det verkliga och centrala problemet när det gäller mellanöstern .
ögonblicket är nu inne , ärade kolleger , att lösa upp en av knutpunkterna när det gäller den globala jämvikten .
ögonblicket är nu inne för israel att hålla sina gamla löften och slutgiltigt dra sig tillbaka från de områden man ockuperat och slutgiltigt och en gång för alla erkänna den palestinska myndigheten , vars återupptagna diplomatiska verksamhet utan tvekan kommer att ha en framtid så länge den befinner sig i yasser arafats erfarna händer .
det är lika viktigt att vi inte förlorar den irakiska frågan ur sikte , en fråga som ingen längre talar om utan man förtränger problemen för miljontals kvinnor , gamla och barn , offer för ett embargo som är lika arrogant som gement .
jag vet inte vad syrien och israel verkligen skulle vilja eller skulle kunna göra , men jag vet att vår institution skulle kunna göra mycket och det är på tiden att vi ägnar oss åt hur människor lever med samma kraft vi som vi ägnar oss åt tändanordningarna till våra lika kalla som vaga och artificiella neonlampor , som kan lysa upp ett hus , men verkligen inte världen under tredje millenniet .
herr talman ! den israeliska författaren , amos oz , beskrev nyligen mycket träffande det kyliga förhandlingsklimatet mellan israel och syrien .
oz hade fått intrycket att syrierna ansåg att de i utbyte för golanhöjden endast behövde faxa ett mottagningsbevis till israelerna .
den tanken av oz dyker också upp i den israeliska pressen .
den återger kontrasten mellan premiärminister baraks personliga fredsansträngningar och den reserverade hållningen , den rent av fysiska frånvaron , hos damaskus starke man , president assad , vid förhandlingsbordet i förenta staterna .
det var väl ändå assad som skulle vara baraks samtalspartner och inte hans utrikesminister .
när det gäller minister farouk al-sharas beteende i shepherdstown är israelerna mycket upprörda .
hans hållning gentemot premiärminister ehud barak var rent ut förnedrande .
vadan denna uppmärksamhet för elementära diplomatiska umgängesformer i en seg territoriell förhandlingsprocess ?
jo , syrierna förstör bara för sig själva .
när allt kommer omkring är det de israeliska väljarna som skall uttala sig om huruvida golanhöjderna skall lämnas tillbaka .
i alla resolutioner som lagts fram uttalas en djup önskan om en större europeisk roll i fredsprocessen .
det är dock frågan om bryssel kan skaffa fram de miljarder dollar som de israeliska och syriska myndigheterna är ute efter hos sin fredsbeskyddare , förenta staterna . då talar vi ändå inte om de tunga , lika dyra säkerhetsgarantierna om israel drar sig tillbaka från golan .
slutligen en fråga till rådet och kommissionen .
vad är sant i pressens uppgifter om att det portugisiska ordförandeskapet redan utlovat trupper till en fredsbevarande styrka i golan ?
sanningen är att brytningen eller förseningen sine die av de pågående samtalen mellan syrier och israeler inte är en bra nyhet . det är inte heller en bra nyhet att ett nytt bombattentat inträffade i förrgår och 16 personer skadades .
det är tydligt att förenta nationerna för en gång skull inte har lyckats i sina medlingsförsök , och det är faktiskt svårlösta hinder . syrierna försöker än en gång att få golan under sin suveränitet och jurisdiktion och få tillbaks de gränser som gällde före den 4 juni 1967 medan israelerna vill ha gränserna dragna som de var 1923 , eftersom det är bättre för dem .
avbrottet i samtalet mellan syrierna och israelerna är inte den enda förseningen i fredsprocessen i mellanöstern .
just nu har tillämpningen av ramavtalet mellan palestina och israel också hävts .
efter samtalen i förrgår mellan israels premiärminister och palestinas ledare begärde den israeliska premiärministern en två månader lång ajournering från och med den 13 februari , sista dag för verkställandet av ramavtalet om situationen på västbanken och gazaremsan .
vad kan europeiska unionen göra i en sådan här situation ? inte mycket , tyvärr .
vi måste givetvis stödja förhandlingarna ledda av förenta staterna .
vi måste intensifiera våra kontakter . europeiska unionens sändebud , ambassadör moratinos , har inom ramen för europeiska unionens befogenheter utfört sitt uppdrag med stor omsorg och effektivitet .
detta till trots kan vi ana en viss maktlöshet , när de båda förhandlingspartnerna i helgen tar flyget hem till förenta staterna får vi inte förglömma att för varje 100 dollar som spenderas i fredsprocessen kommer 60 från europeiska unionen .
när vi dessutom beaktar att nästa möte kommer att hållas i moskva , så blir europeiska unionens närvaro något patetisk .
inför det portugisiska ordförandeskapet insisterar jag på en mera central roll , det är dags för europeiska unionen att ta över och bli mera delaktig .
jag hoppas att nästa besök i regionen av europaparlamentets talman , samt av de interparlamentariska delegationerna och deras ordförande , tillåter oss att inleda en mera initiativrik etapp där europeiska unionen tydligare kan delta i denna komplicerade och svåra fredsprocess .
herr talman , herr rådsordförande , kommissionär patten ! jag vill tacka för era redogörelser , särskilt gäller det kommissionär patten vars analys jag helt och fullt delar .
jag kommer av den anledningen ej att upprepa något av vad han sagt . i stället vill jag göra tre kommentarer som kommissionär patten måhända har samma syn på men som han av olika skäl inte kan formulera lika öppet som en ledamot kan göra .
det första är att jag tror att vi har anledning att glädja oss över det avtal som finns mellan israel och den palestinska myndigheten för självbestämmande .
nu finns det dock tillräckligt med avtal : oslo , wye plantation , sharm-el-sheik .
det räcker så , nu måste de uppfyllas också .
på den punkten delar jag emellertid min kollega salafrancas skepsis när han säger att det kom dåliga nyheter från israel , närmare bestämt att även detta senaste avtal inte kommer att kunna uppfyllas i tid .
den andra punkten gäller återupptagandet av förhandlingarna mellan syrien och israel .
detta är , menar jag , en högst glädjande nyhet .
men denna vecka har vi också fått höra att barak inte reser till washington och att förhandlingarna därmed inte kan fortsättas .
jag vill klart och tydligt slå fast att om golanhöjderna lämnas tillbaka till syrien så är problemet löst i denna region .
gällande frågan om folkomröstning som berörts av flera kolleger : vi måste nu fråga oss om man verkligen alltid måste hålla folkomröstning för att kunna uppfylla förpliktelser ur internationell rätt och folkrätten .
i tyskland skulle man förmodligen glädja sig mycket om vi sade att vi genomför en folkomröstning för betalningen till europeiska unionen ; men vi gör det oberoende av huruvida det tyska folket är villigt att betala .
det skulle vara en likartad situation .
min tredje och sista punkt gäller europeiska unionens roll .
här vill jag verkligen framhålla den enastående roll som det särskilda sändebudet moratinos har spelat i regionen , samt även det vi åstadkommit i form av finansiering , kommissionär patten .
ni skall veta att ni alltid kan få stöd för ert förslag i detta parlament . vi kommer att finnas där när det skall finansieras .
vi bör dock också spela en politisk roll , som ju moratinos inte kan göra helt själv i denna region . rådsordförandeskapet måste då aktiveras , mister gasp måste då ta sig till regionen , och vi måste själva bjuda in förespråkarna för fredsprocessen , på samma sätt som ryssarna gjort .
då har vi tagit det ansvar som motsvarar vårt engagemang och bidrag .
herr talman , kommissionär patten , kära kolleger !
de senaste fredsförhandlingarna som inletts i förenta staterna mellan israel och syrien är en vändpunkt i mellanösterns historia , en vändpunkt som man väntat på i femtio år nu och som uppenbarligen är svår att förhandla om .
det blir inget möte i dag i shepherdstown , men vi skall hoppas , såsom kommissionär patten nyss sade , att detta uppskjutande av förhandlingarna på grund av de senaste kraven från syrien , bara är en incident på vägen mot ett fredsavtal som kan ändra hela mellanösterns utseende .
det är vad vår resolution uttrycker : en förhoppning om ett rimligt och rättvist avtal , grundat på respekt för de suveräna staterna och rätten att leva i säkerhet inom säkra och erkända gränser .
alla utländska trupper , inbegripet de syriska , måste alltså lämna libanon , i enlighet med resolution 520 från förenta nationernas säkerhetsråd .
kan vi hoppas på att vi i juli 2000 - det datum som ehud barak lovat - fått uppleva en israelisk reträtt ur södra libanon ?
kan unionen hoppas på ett dubbelt fredsavtal mellan israel och dess grannar i norr ?
vi tror det . vi vill tro det .
aldrig har parternas beslutsamhet varit starkare .
jag skulle också vilja betona en punkt som förefaller mig grundläggande : balansen som måste känneteckna vårt europeiska budskap , en politisk balans mellan dem som deltar i förhandlingarna naturligtvis , men också balans mellan befolkningarna .
efter attentatet mot hadera i måndags måste vi upprepa vårt fördömande av varje form av terrorism .
och apropå balans , eller obalans snarare i detta sammanhang , skulle jag vilja lägga till hur beklagligt det är att återigen tvingas konstatera vilken svag politisk roll europa spelar när det gäller att lösa konflikten .
vid lunchtid i dag tog rådets ordförande gama upp europas ekonomiska och handelsmässiga stöd till regionen .
man måste trots allt konstatera att inledandet av fredsprocessen för närvarande i huvudsak är washingtons verk .
syrierna har , liksom andra arabiska länder före dem , valt ut amerikanerna för att beskydda förhandlingarna .
det är också det val den hebreiska staten gjort där europa , det är ett faktum och inte någon bedömning , lider av en partisk offentlig bild .
det är alltså rätt tillfälle att på nytt säga till kommissionär patten , till solana och till moratinos , att vi verkligen räknar med deras ansträngningar för att den europeiska rösten skall höras , i strävan efter en fredlig lösning av konflikten .
och även om det är svårt för europa att tala med en röst om fredsprocessen kan , och måste vi , ändå tala om den i samma anda av förtroende och solidaritet .
nästa punkt på föredragningslistan är muntliga frågor till rådet ( b5-0040 / 99 ) och till kommissionen ( b5-0041 / 99 ) från utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikes frågor om årsrapporten 1999 och om området frihet , säkerhet och rättvisa ( artikel 39 i maastrichtfördraget ) .
mina damer och herrar , ärade rådsmedlemmar ! för det första , utan att gå in på någon tävling om känslor med ministrarna , vill jag säga att jag inte känner sinnesrörelse , jag känner mig förvirrad av att i ordförandeskapet för första gången ha två personliga vänner och jag hoppas att detta faktum inte kommer att förändra maktdelningen , som är viktig för vår union .
sedan skulle jag vilja gratulera ledamoten anna terrón till att ha tagit upp den fråga som gett upphov till den första debatten i år under denna mandatperiod om skapandet av ett område med frihet , säkerhet och rättvisa , samt tacka alla ledamöter som i de olika utskotten har deltagit aktivt i förberedandet av denna debatt , liksom företrädarna för de nationella parlamenten och det civila samhället .
jag vill i detta första inlägg ge parlamentet kommissionens syn på det mest betydelsefulla som hände under år 1999 .
jag tycker att jag med övertygelse , men också med tillfredsställelse , kan säga att år 1999 var en vändpunkt och ett befästande av unionen i frågorna om frihet , säkerhet och rättvisa .
det har redan sagts här att amsterdamfördraget trädde i kraft i maj , och detta parlament ansåg att den mest långtgående nyheten i detta fördrag var erkännandet av att det var nödvändigt att skapa ett område med frihet , säkerhet och rättvisa .
detta utgör samtidigt ett kvalitativt mycket viktigt hopp framåt och ett logiskt och oumbärligt steg i unionens utveckling , efter skapandet av den inre marknaden , införandet av den gemensamma valutan och lanserandet av en gemensam utrikes- och säkerhetspolitik .
detta projekt är , mer än ett institutionsprojekt , ett projekt för medborgarna i vår gemensamma union .
därför måste alla medborgare i unionen få en verkligt fri rörlighet , och vi måste erkänna att denna bara är meningsfull om den genomförs i ett säkert sammanhang , med stabil grund i ett effektivt rättsligt system som alla har tillgång till under enkla och lika förutsättningar , och som medborgarna kan lita på .
unionens ansträngningar att förverkliga ett område med frihet , säkerhet och rättvisa befästes i tammerfors .
jag skulle vilja understryka det starka politiska budskap som europeiska rådet gav , där det framhöll den betydelse stats- och regeringscheferna lade vid ett viktigt förslag , liksom vid antalet politiska riktlinjer och prioriteringar som kommer att göra detta område verkligt , enligt en progressiv strategi , inom ett femårigt perspektiv och detta område har framför allt tre beståndsdelar : frihet , säkerhet och rättvisa .
år 1999 präglades också av det tyska ordförandeskapets initiativ att utarbeta en stadga om grundläggande rättigheter i unionen .
i europeiska unionens nuvarande utvecklingsfas , anser jag att det vore lämpligt att samla de gällande grundläggande rättigheterna på unionsnivå i en stadga , för att göra dem mer synliga och tillgängliga för alla medborgare .
som jag redan har sagt flera gånger så är jag för , och kommissionen är för , att utarbeta en stadga som , grundad på en dynamisk process , återspeglar medlemsstaternas gemensamma konstitutionella traditioner och de allmänna principerna i gemenskapsrätten , och inte bara reducerar dem till en formulering med minsta gemensamma nämnare .
som företrädare för kommissionen kommer jag att vaka över att stadgan och dess åtgärder befäster en union , som grundas på en rad grundläggande rättigheter som är en del av europas gemensamma arv .
bara så kan vi bidra till att legitimera utvidgningsprojektet av unionen i alla europeiska medborgares ögon , en utvidgning som grundas på respekten för rättigheter och friheter , en garanti för människors och egendoms säkerhet och med ett effektivt rättsligt skydd , det vill säga , en union som är grundad på politiska värden som de nuvarande demokratierna bygger på .
jag tänker inte utelämna att 1999 också var det år då mandatperioden 1999-2004 inleddes i europaparlamentet och den nya kommissionen tillträde och därmed en kommissionär med exklusivt ansvar för det rättsliga och inrikes området .
förutom dessa händelser , skulle jag vilja påminna parlamentet om några saker som antogs under år 1999 .
kommissionen lade fram ett förslag till förordning i fråga om invandring , gränser och asyl , för skapandet av databasen &quot; eurodac &quot; , förslaget till direktiv om villkoren för tredjelandsmedborgares inresa och vistelse i unionens medlemsstater för att återsamla familjer , inom ramen för en bestämd integrationspolitik av dem som vistas legalt i unionen .
vi satte i gång en debatt om ett meddelande om gemensamma förfaranden angående asyl och en rekommendation till beslut som bemyndigar kommissionen att förhandla om ett avtal med island och norge om en utsträckning av de bestämmelser som europeiska unionens medlemsstater tillämpar enligt dublinkonventionen till dessa båda länder .
kommissionen bidrog aktivt till arbetet i högnivågruppen om asyl och invandring och slutligen , i december , lade den fram ett förslag till skapandet av europeiska flyktingfonden .
på området för rättsligt samarbete lade kommissionen fram förslag till förordningar för att göra vissa konventioner till gemenskapsfrågor : om rättsligt samarbete och verkställighet av domar av civil eller kommersiell natur , ( bryssel-i ) ; en annan , angående erkännande och verkställighet av domar i äktenskapsmål ( bryssel-ii ) och ännu en annan , delgivning i medlemsstaterna av handlingar i mål och ärenden av civil eller kommersiell natur .
vi lade också 1999 fram ett meddelande om brottsoffer i unionen och inledde därigenom en diskussion som i tammerfors tog ett steg framåt och som innehåller krav på minimibestämmelser om skydd för brottsoffer , speciellt tillgång till rättslig hjälp och rätt till ersättning för skador , inklusive rättsliga kostnader .
jag vill också nämna förslaget till beslut om åtgärder för att bekämpa bedrägeri och förfalskning som rör andra betalningsmedel än kontanter .
inom ramen för unionens lagstiftning om ekonomisk brottslighet , lade kommissionen fram ett förslag till revidering av direktivet om penningtvätt .
vi deltog 1999 i starten av europol , och från kommissionen hoppas vi uppriktigt , särskilt efter vad det portugisiska ordförandeskapet sade här i dag , att den nya perioden för rättsliga och inrikes frågor , och de påbörjade diskussionerna om att införa nya befogenheter för europol i amsterdamfördraget , också skall följas av en diskussion om demokratisk kontroll och förbindelserna mellan europol och behöriga rättslig instans , nämligen eurojust .
kommissionen lade 1999 även fram sitt bidrag till en europeisk handlingsplan för narkotikabekämpning , vilken ligger till grund för den strategi som godkändes av europeiska rådet i helsingfors .
denna åtgärdslista , som inte är uttömd , har bidragit till att jag i dag , inför rådets ordförandeskap och ledamöterna , med stor övertygelse kan säga att , om 1999 var ett år som befäste unionens verksamhet inom detta grundläggande område så hoppas jag också att 1999 innebär början på en ny period , en strävan att skynda på skapandet av ett område med frihet , säkerhet och rättvisa .
därför kommer år 2000 utan tvivel att bli ett år för att pröva hur de europeiska institutionerna klarar att möta medborgarnas krav om fri rörlighet , i respekten för rättigheter och i garantier för säkerhet och stabilitet , genom ett adekvat rättsligt skydd .
vi kan också säga att år 2000 för rådet , parlamentet och kommissionen kommer att vara ett prövoår för den politiska viljan att ta amsterdam på allvar och lägga grunden för en utvidgad politisk union under nästa decennium .
som jag har sagt är kommissionen medveten om sin del av ansvaret och i detta sammanhang har den snart avslutat ett första utkast till förslag till resultatöversikt , en scoreboard , där alla institutioner och andra berörda delar kan börja utvärdera de framsteg som skett genom införandet av nödvändiga åtgärder och uppfyllandet av de tidsfrister som fastställts i amsterdamfördraget , handlingsplanen från wien och slutsatserna från tammerfors .
denna resultatöversikt kommer inte bara att vara ett instrument för programplanering av lagstiftning utan också , och framför allt , ett instrument för att stärka alla europeiska institutioners öppenhet och ansvar inför medborgarna .
detta därför att det är för medborgarna som vi utvecklar ett område med frihet , säkerhet och rättvisa .
framstegen beror inte på kommissionen , inte på rådet , inte ens på europaparlamentet , utan på de europeiska institutionerna i helhet och på medlemsstaterna själva , då vissa uppgifter på resultatöversikten , vilket redan har sagts här , anförtros medlemsstaterna enligt subsidiaritetsprincipen .
de närmaste veckorna kommer jag att genomföra en rundresa i huvudstäderna för att lyssna på ministrarna för rättsliga och inrikes frågor .
jag räknar med att debattera projektet med resultatöversikt med europaparlamentet och med det civila samhället .
vi räknar med att efter dessa konsultationer lägga fram slutversionen inför rådet för justitie- och inrikesministrar , under det portugisiska ordförandeskapet .
min avsikt är att denna resultatöversikt skall bli ett instrument för politisk och strategisk inriktning för alla institutioner men också ett instrument för opinionsundersökningar .
därför inser jag - och det är en utmaning som jag tror att vi alla ställs inför - , att utveckla en kommunikationsstrategi som kan göra det mervärde som unionen innebär för allmänheten i dess dagliga liv , tillgängligt och begripligt i dessa viktiga områden för medborgarna , i respekten för lagligheten och i grunden själva demokratin .
förutom resultatöversikten skulle jag vilja nämna att kommissionen räknar med att under år 2000 lägga fram följande initiativ - och jag skulle här vilja understryka att jag gratulerar till att det portugisiska ordförandeskapet betraktar utvecklingen av detta område som en av sina prioriteringar i arbetsprogrammet .
jag hoppas att det blir möjligt , under det portugisiska ordförandeskapet , att tydligt utveckla en interinstitutionell samarbetsanda , vilket också är det politiska budskapet från tammerfors , och att denna interinstitutionella samarbetsanda följs upp av de efterföljande ordförandeskapen .
när det gäller invandring och asyl , räknar kommissionen med att kunna lägga fram förslag till utformningen av ett gemenskapsinstrument för tillfälligt skydd av flyktingar ; inleda analysen av kriterier och villkor för att förbättra genomförandet av dublinkonventionen och ett övervägande att förändra dess rättsliga grund i enlighet med amsterdamfördraget ; fortsätta debatten utifrån det meddelande som redan har spridits om bestämmelser som leder till ett gemensamt asylförfarande i hela unionen ; och lägga fram lagstiftningsförslag om att bevilja uppehållstillstånd till de offer för människohandel som samarbetar med rättsväsendet mot nätverken för människohandel .
jag räknar också med att kunna bidra till ett klargörande av handlingsplanernas roll inom arbetet i högnivågruppen om asyl och invandring och gå vidare med antagandet av gemenskapsavtal för återinresa , genom att införa klausuler för detta ändamål .
i en central fråga angående den fria rörligheten såsom resa över de yttre gränserna i medlemsstaterna kommer jag under de närmaste dagarna att lägga fram ett förslag till förordning som förnyar listan över tredje land vars nationaliteter måste ha visering för att kunna passera de yttre gränserna .
inom det rättsliga samarbetet hoppas jag innerligt att det , förutom ett initiativ om lagen som är tillämplig på förpliktelser ej angivna i kontrakt blir möjligt att lägga fram ett förslag till minimibestämmelser som garanterar en lämplig nivå av rättshjälp över hela unionen vid gränsprocesserna .
jag räknar också med att kunna fortsätta arbeta med nya gemensamma processregler specifikt för att förenkla och påskynda av gränsöverskridande rättsliga processer i mindre fall gällande handel och konsumenter , matpensioner och ej besvarade åtal .
i uppföljningen av slutsatserna från tammerfors och helsingfors kommer kommissionen att lägga fram sitt bidrag till definitionen av en unionens strategi för att förebygga och bekämpa den organiserade brottsligheten .
vi kommer att organisera och stödja åtgärder och särskilt debatten om behovet att utarbeta ett lagstiftningsprogram för genomförande av principen om ömsesidigt erkännande av domar i straffrätten .
kommissionen räknar också med att lägga fram specifika åtgärder för förebyggande av brottslighet för att utveckla utbytet av den bästa praxisen på området , speciellt förebyggande av brottslighet i städerna och ungdomsbrottslighet , och lägga fram en rättslig grund för ett program , finansierat av gemenskapen .
kommissionen kommer också att bidra till ordförandeskapets arbete för att klargöra den rättsliga ramen och den administrativa polisiära och rättsliga samarbetsramen för att bekämpa penningtvätt , i ett perspektiv som i hög grad överskrider gränserna mellan pelarna .
kommissionen kommer att uppfylla det ansvar den fick i tammerfors för att lägga fram förslag till antagande av gemensamma definitioner , åtal och sanktioner mot människohandel och ekonomiskt utnyttjande av invandrare och sexuellt utnyttjande av kvinnor och barn , med särskild tonvikt lagd på kampen mot användande av de nya kommunikationsmedlen , främst internet , för spridning av barnpornografi .
vi förbereder också ett meddelande för att diskutera medlen för att skapa ett samhälle med säkrare information och kunskap och för att kunna bekämpa datorbrottslighet .
år 2000 innebär också inledningen av tillämpningen av den europeiska strategin mot narkotika för perioden 2000-2004 .
kommissionen kommer på detta område och i samarbete med det portugisiska ordförandeskapet och europaparlamentet , att ge allt sitt stöd till den interinstitutionella konferensen i februari om narkotikaproblematiken .
beträffande schengen skulle jag , utan att nu gå in på rådets behörighetsområde , och särskilt när det gäller integreringen av schengenregelverket inom gemenskapsramen , vilja understryka att kommissionen , i den aktuella frågan om återupprättandet av gränskontroll , än en gång upprepar sin beredskap att fördjupa formerna för en bättre kontroll av tillämpningen av artikel 2.2 i schengenkonventionen , så att den blir mer tvingande .
återinrättandet av viss intern gränskontroll nyligen får mig att dra slutsatsen att det är nödvändigt att göra en detaljanalys av förutsättningarna för att anta ett lagstiftningsinstrument grundat på artikel 62 i fördraget .
så som betonades i tammerfors , och med tanke på förberedelserna av europeiska rådet i feira , i juni 2000 , måste vi sammanfatta innebörden av den nya externa dimensionen i de inrikes och rättsliga frågorna med perspektiv på ett antagande av politiska strategier mellan pelarna för att förstärka sammanhållningen i unionens inrikes- och utrikespolitiska förbindelser för att bidra till att befästa unionen i världen .
jag vill emellertid understryka att alla dessa åtgärder givetvis måste ske med hänsyn till de principer som beslutats vid europeiska rådet i helsingfors i förhållande till ansökarländerna , så att dessa ansökarländer samarbetar och så snart som möjligt knyts till projektet att skapa ett område med frihet , säkerhet och rättvisa .
det är för övrigt viktigt att komma ihåg att förhandlingarna om rättsliga och inrikes frågor inleds år 2000 med den första gruppen ansökarländer och jag hoppas att vi skall kunna göra stora framsteg i förberedelserna av de förhandlingsärenden angående den andra gruppen som i helsingfors godkändes för anslutning .
slutligen skulle jag vilja säga att kommissionen försöker vara i en pole position i presentationen av förslag för att kunna följa upp genomförandet av amsterdamfördraget .
jag hoppas att kommissionen och rådet kommer fram till ett avtal om delat ansvar i utövandet av initiativrätten och ledningen av själva lagstiftningsprocessen .
som jag sade till parlamentet , den uppgift vi har framför oss är enorm och ambitiös , kommissionen behöver vara utrustad med nödvändiga mänskliga resurser för att kunna möta denna utmaning och hoppas få parlamentets stöd , och varför inte rådets , för att garantera dessa resurser och mål , så att skapandet av ett område med frihet , säkerhet och rättvisa i unionen blir verklighet så snart som möjligt och på så sätt kan vi alla bidra , i en anda av interinstitutionellt samarbete , för att genomföra detta projekt , vilket utan tvivel är &quot; kronjuvelen &quot; i amsterdamfördraget .
efter att denna församling under 40 år ägnat sig huvudsakligen åt att etablera en gemensam inre marknad har vi nu en ny stor uppgift i att skapa ett område av frihet , säkerhet och rätt . det är en uppgift som vi emellertid endast kommer att kunna lösa framgångsrikt om alla unionens institutioner arbetar gemensamt med ömsesidig respekt mot det ambitiösa målet , under beaktande av respektive befogenhetsområden .
kommissionär vitorino , medan jag vill beteckna samarbetet med er som harmoniskt och fruktbart så har jag ofta saknat ord för att beskriva det uppträdande som rådet visat prov på i förbindelserna med oss .
det har verkat - som kollegan schulz en gång träffande sagt i utskottet - som om rådet under området av frihet , säkerhet och rätt tänkt sig ett område för egen oansvarighet , för säkerhet att inför parlamentet och rätten göra och låta ske enligt eget godtycke .
herr minister gomes , jag har förstås uppfattat era redogörelser om detta . följaktligen hoppas jag på en tydlig förbättring i samarbetet under det portugisiska rådsordförandeskapet .
jag vill lyfta fram tre punkter vilka för oss medlemmar i europeiska folkpartiets grupp måste vara tyngdpunkter i skapandet av ett sådant område .
för det första : uppbyggandet av en gemensam asylrätt och en fördelning av de bördor som uppkommer i samband med mottagande av flyktingar .
först måste rådet äntligen tillse att eurodac blir utfärdat för att skapa en grundförutsättning för fördelning av asylsökandena .
vad beträffar en asylrätt som gäller över hela europa har förvisso ett par ansatser blivit synliga genom wien och tammerfors .
dessa ansatser visar emellertid dessvärre snarare på de svårigheter som finns i stället för att komma med lösningsförslag .
företrädarna i rådet uppmanas därför att blicka ut över sina egna nationella murar och skapa ett enhetligt asylförfarande för hela unionen .
det kan heller inte vara riktigt att några få hjälpvilliga medlemsländer skall tvingas bära hela bördan av flyktingeländet på vår kontinent .
en överenskommelse om en fördelning av bördorna måste av den anledningen ha högsta prioritet .
för det andra : utbyggnaden av ett alleuropeiskt bekämpande av den organiserade brottsligheten , bland annat via europol och eurojust .
det planerade inrättandet av eurojust framstår för oss som ett viktigt framsteg från tammerfors som nu måste genomföras snarast .
vi välkomnar det faktum att europol till slut har kunnat påbörja sitt arbete .
rådet får dock ej bortse från att det för att effektivisera brottsbekämpningen inte räcker med den i tammerfors beslutade fördelningen av europols uppgifter , utan att det måste ingå såväl en personell förstärkning som en uppgiftsfördelning ända ned till den operativa nivån .
det är inte så att vi ropar efter ökad kontroll och mer kontroll över själva europol ; för oss gäller här snarare talesättet : &quot; mindre är ibland mer ! &quot;
om en huvuddel av europols medarbetare för närvarande framför allt är sysselsatta med att kontrollera sig själva i datasäkerhetsrättsligt hänseende varvid man inhämtar undersökningar från 15 olika nationella parlament är detta mycket kontroll , men en ineffektiv kontroll .
vi vill ha mindre virrvarr i kontrollen men ökad parlamentarisk kontroll genom europaparlamentet , och detta utan att europols arbete skall hindras .
samtidigt stöder vi inrättandet av en europeisk polisakademi , vilket föreslagits i tammerfors , såsom ett steg i rätt riktning .
för det tredje : utvidgningen av parlamentets rättigheter i detta sammanhang .
om det bara blir diplomater och byråkrater som bestämmer över inrättandet av en anordning som medger unionen att även ingripa i de grundläggande fri- och rättigheterna för unionens medborgare , medan de valda företrädarna i europa inte kan annat än bara följa utvecklingen som kaniner gör med ormens rörelser , så kommer denna anordning aldrig att accepteras av medborgarna .
det är därför på tiden att parlamentet härvidlag tillerkänns medbeslutanderätt och - som redan sagts - att principen om demokratisk kontroll stärks .
vi vill ha ett område av frihet , säkerhet och rätt för medborgarna i europa och inte mot dem .
jag välkomnar varmt det faktum att det portugisiska ordförandeskapet sätter rättsliga och inrikes frågor högt , om inte högst , på prioriteringslistan .
jag blev också glad att höra kommissionär pattens kommentarer i förmiddags om en fond för snabba åtgärder vid säkerhetskriser .
kanske detta kan få slut på skandaler som misslyckandet med att sätta in den utlovade polisstyrkan i kosovo .
låt mig bara betona tre områden bland många där vi behöver se snabba framsteg .
det första rör asyl .
det är nödvändigt att upprätta ett gemensamt europeiskt system , men det skall grundas på rättvisa , fullständig respekt för genèvekonventionen och anständiga mottagningsförhållanden , inklusive ett slut på de rutinmässiga kvarhållandena .
ett asylbeslut bör kunna fattas inom några månader - inte inom några år .
det andra området rör frihet : frihet att flytta och bosätta sig var man vill inom unionen ; informationsfrihet ; frihet att rösta på alla som har ett europeiskt medborgarskap - och detta omfattar inte bara medborgare i medlemsstaterna , utan även medborgare från tredje land .
låt våra medborgare få veta att vår gemensamma politik rörande rättsliga och inrikes frågor handlar om frihet , inte bara om förtryck .
det sista området jag vill nämna handlar om konvergering av civil- och straffrättsliga system .
euroskeptikerna hävdar att detta är ett hot mot suveräniteten , slutet för nationalstaten , osv. men fallet som rör den misstänkte som var efterlyst för utfrågning i samband med morden på tre kvinnor i frankrike , inklusive den brittiska studentskan isabel peake , som blev avslängd från ett tåg , visar varför vi behöver ett ömsesidigt erkännande .
mannen som arresterades och släpptes i madrid , har nu blivit utlämnad efter att ha suttit arresterad i lissabon .
vad euroskeptikerna än säger ligger det i allas vårt intresse att det sker ett samarbete kring sådana frågor .
sammanfattningsvis , som redan nämnts , är det nödvändigt - och jag hoppas att detta tas upp på regeringskonferensen - att det ändras till medbeslutandeförfarandet inom dessa områden , med demokratisk och rättslig granskning .
herr talman , angående år 1999 kan jag bara säga följande helt kort : efter den finska kylan är portugals solsken hjärtligt välkommet .
jag hoppas att det också går bra .
en för europa viktig händelse under 1999 när det gäller området av frihet , säkerhet och rättvisa var helt säkert toppmötet i tammerfors .
men fortfarande kvarstår åtskilliga frågor att besvara .
många svar väntar vi ännu på .
dock efter tammerfors har vi fått en obalans mellan de positiva åtgärder som faktiskt vidtogs och rena avsiktsförklaringar .
det återstår fortfarande att besluta om medborgarskapsregleringen samt om integrationen av människor från tredje land .
å andra sidan har man nu tagit initiativ till högst konkreta åtgärder på temat säkerhet .
framtagandet av en stadga med grundläggande fri- och rättigheter torde bli ett av de stora projekten i den nära framtiden .
när jag tänker på de människor som för närvarande ej är unionsmedborgare känns det dock svårt att förutsäga hur denna stadga kommer att se ut rent innehållsmässigt och vilken utformning i rättslig mening förverkligandet av den kommer att få .
europolavtalet har nu officiellt trätt i kraft .
vid mötet i tammerfors siktade man på att också fördela de operativa befogenheterna .
men vi kräver alltjämt en revidering av avtalet , vilket syftar till att åstadkomma förbättrade parlamentariska och rättsliga kontrollmöjligheter .
också vad gäller eurodac bör avtalet ställas under kritisk belysning .
parlamentet har modifierat fördragstexten .
det måste garanteras att rådet går på samma linje som parlamentet .
vad gäller övriga ämnen har det tyvärr ännu inte tagits några initiativ . vi väntar för ögonblicket på det .
europa såsom ett område av frihet , säkerhet och rättvisa är fortfarande en anordning utan klar reglering på centrala områden .
vi är dock skyldiga de europeiska medborgarna detta .
efter att ha hört inrikesministern och justitieministern tala är jag numera optimistisk . jag utgår ifrån att vi kommer att lyckas med detta under de kommande sex månaderna .
jag tror att den muntliga frågan från terrón i cusí är intressant så till vida att den är ett tramp i klaveret , för sex månader efter att vårt nya parlament inrättats måste vi kunna ge ett starkt politiskt budskap till europas medborgare .
jag tror att det portugisiska ordförandeskapet positivt kan bidra till det .
vi känner i dag alla till de ofantliga förväntningarna från våra landsmän när det gäller frihet , säkerhet och rättvisa , bl.a. på det sociala området .
men deras brist på intresse , deras distans och ibland t.o.m. avsky för politiken tvingar oss att vidta konkreta åtgärder mot svårigheterna .
det är ett oeftergivligt villkor för att de på nytt skall komma överens med politiken .
för att europa skall bli en symbol för fred och broderskap måste vi bedriva en djärv och generös politik och hjälpa de sämst lottade .
en verklig handlingsplan mot arbetslösheten måste inrättas , för det är utifrån denna farsot som rasism , främlingsfientlighet , nationalism och den rasistiska extremhögern frodas .
bland de sämst lottade , och det är viktigt att jag nämner den punkten , har vi invandrarna och flyktingarna .
villkoren för att praktiskt taget systematiskt kvarhålla och kriminalisera asylsökande är inte längre godtagbara .
alla asylsökande måste få rätt att höras rättvist och ha rätt till suspensiv talan .
jag blev av en tillfällighet vittne till en scen med sällsynt våld i förra veckan på roissys flygplats , där två unga kvinnor , säkerligen illegala invandrare , återfördes till conakry .
de behandlades som de värsta brottslingar .
de var nakna , släpades i håret över golvet och omringades av en hord kravallpoliser .
det portugisiska ordförandeskapet måste få ett stopp på detta slag av barbariska vanor .
vår roll är i stället att åtfölja , garantera , hjälpa dem som flyr från diktaturer .
kommissionen föreslog att en europeisk fond för flyktingar skulle inrättas . parlamentet är mycket positivt till det .
i stället för att komma med undanflykter när det gäller den budget som beviljats fonden tror jag ni kan fatta beslutet att inrätta den .
ordförandeskapet och rådet kan konkretisera det som förkastats som obegripligt i tammerfors , även om tammerfors utgjorde en viktig grund .
på samma sätt kan vi inte nöja oss med att konstatera att de främlingsfientliga strömningarna ökar i europa och att man banaliserar diskriminering , utan att vidta omfattande åtgärder .
det krävs harmonisering av lagstiftningen mot rasism .
vilken inriktning vill ni ge artikel 13 i fördraget ?
vad tänker ni göra för att främja lika lön för män och kvinnor ?
hur tänker ni arbeta för att utrota homofobin , rasismen och sexismen ?
vi måste använda de bästa tillämpningarna från varje land i unionen .
när sex europeiska länder beviljar rösträtt kan er president tillåta sig att utvidga denna rösträtt och valbarhet i de kommunala och europeiska valen till samtliga medborgare från länder utanför unionen , som sedan fem år bor på europeiskt territorium .
att ge de personer som inte har några identitetshandlingar uppehållstillstånd i vissa länder , däribland ert , måste bli ett exempel för de övriga , för denna grupp utan identitetshandlingar består i dag av sköra människor som befinner sig i händerna på utsugare och som utnyttjas som arbetskraft , vilket gör dem till den moderna tidens slavar .
rent allmänt måste detta ordförandeskap inleda förändringar när det gäller uppträdande och förhållanden bland våra landsmän tillsammans med minoriteter och invandrare .
immigrationen är alltför ofta synonym med osäkerhet och våld och rent repressiva lösningar .
hur skall ni få våra landsmän att förstå att immigrationen i dag , liksom alltid , är en källa till social och kulturell rikedom , vars roll är och förblir nödvändig i vår demografiska miljö .
vilka åtgärder avser ni att vidta för att uppvärdera invandrarnas plats i samhället och garantera ett verkligt skydd för asylsökande ?
herr talman ! det råder stor brist på öppenhet inom området säkerhet , frihet och rättvisa .
europeiska unionen är en ekonomisk jätte , men vi har inte rätt att spela ofelbara när det gäller vår behandling av flyktingar .
nivån på rasismen i vårt samhälle är skrämmande .
under flera generationer skickade irland iväg sina söner och döttrar till säkra platser över hela världen , men nu när den keltiska tigern skapar ett välstånd som är större än vad vi förväntat oss , visar vi ett mycket fult drag i vår karaktär .
rasismen i irland är endemisk .
det var en ganska stor chock för våra politiska ledare när de förstod att vi nu måste ta en del av de flyktingar som under en lång tidsperiod rest till europeiska unionen .
vi har kommit efter när det gäller att ta itu med denna fråga och regeringen gör sitt yttersta för att hinna ikapp .
viljan finns , men rädslan dröjer sig kvar ; och för att dämpa denna rädsla måste vi hitta ett politiskt och religiöst ledarskap , inte bara i irland utan över hela europeiska unionen .
herr talman ! vi kan notera att det urskuldande och försiktiga ordförandeskap som under de senaste månaderna har förhindrat en debatt som den vi faktiskt har lyckats genomföra i dag , har upphört .
jag instämmer till fullo i det som mina kolleger von boetticher och schulz sade och anser det vara helt rätt att europaparlamentet och domstolen måste engagera sig mer i området frihet , säkerhet och rättvisa utan att behöva avstå från sina egna befogenheter .
men just för att vi inte skall behöva upprepa det spektakel som var sjätte månad urskillningslöst drabbar rådets ordförande , borde kanske detta parlament ha modet att ta ett kraftfullt politiskt initiativ så att nästa regeringskonferens beslutar att genast utvidga medbeslutandet i stället för att vänta i ytterligare fem år .
de två likalydande frågorna som behandlas , bärs fram av ett mantra som numera mer och mer förvandlar politik till en slags ideologi - välklingande , men fördärvlig .
och våra dagars eu-mantra heter ofsr - område för frihet , säkerhet och rättvisa .
bakom detta ligger en annan ambition hos kommissionen , rådet och det överväldigande flertalet i denna församling , dvs. att införa ett sådant område .
och vem stöder då inte säkerhet , frihet och rättvisa ?
problemet är bara att det inte är något som eu kan införa genom lagstiftning och andra övernationella åtgärder .
frihet , säkerhet och rättvisa är ett samhälles rotsystem . det är en återspegling av varje samhälles historia , dess sociala erfarenheter och politiska utveckling .
det är inte något som eu kan införa utan att samhället lider skada .
men det är just här vi hittar det faktiskt rationella i mantrat om säkerhet , frihet och rättvisa .
uppgiften är inte att säkerställa rättvisa för medborgarna .
det sker redan genom de nationella rättssystemen .
uppgiften är att överföra viktiga delar av samhällets straffrätt , kriminalpolitik och rättskipning till eu : s institutioner .
det handlar om en förstärkt integration som t.o.m. i en bedräglig förpackning innehåller förstärkt repression och kontroll .
tänk bara på alla åtgärder kring fästning europa , schengen , eurodac osv. varje demokrat hittar två nyckelproblem .
för det första är de planerade åtgärderna helt orealistiska .
hur föreställer man sig att eu : s institutioner , som redan lider under en tung arbetsbörda , skall kunna genomföra dessa ambitiösa projekt ?
tänk på de senaste årens mördande kritik av kommissionens brist på anständighet , etik och ansvar .
det kommer ju också till direkt uttryck i frågan .
för det andra är projekten belastande - ja , lemlästande - för de nationella demokratierna .
så länge som eu sysslade med den inre marknaden angrep man bara kroppen .
nu angriper man själen .
herr talman ! i dag har det nordirländska folket fått bevittna en underlig , ironisk händelse .
kommissionär patten har talat i kammaren och försvarat frihet , säkerhet och rättvisa , och trots detta resulterar den rapport han lagt fram för det brittiska underhuset - vilken har accepterats - i att the royal ulster constabulary och dess reserver försvinner och att nordirländare , både protestanter och katoliker , hamnar i händerna på terrorister .
terroristerna från ira har inte lämnat inte några vapen , vilket inte heller de protestantiska terroristerna har gjort , ändå tvingas polisen in i ett läge där de inte har befogenheter att bekämpa terroristerna .
låt mig ta en titt på siffrorna från den dag avtalet undertecknades .
under 1998 hade vi 55 mord .
under 1999 hade vi sju mord och då räknas inte offren för bomben i omagh med , där 29 dödades och 300 skadades .
mellan 1998 och 1999 överföll och sköt lojalisterna 123 personer , medan republikanerna överföll och sköt 93 personer .
antalet åtal som väcktes mot lojalisterna under 1999 uppgick till 193 och motsvarande siffra för republikanerna var 97 .
sedan januari 2000 har det skett sex överfall med skjutvapen som utförts av lojalisterna och två av republikanerna ; lojalisterna har varit inblandade i sex allvarliga överfall , varav ett resulterade i ytterligare ett mord , samtidigt som republikanerna varit inblandade i fem allvarliga överfall .
herr talman ! man måste komma till rätta med situationen - detta kan inte fortsätta .
amsterdamfördraget har visat sig vara ett viktigt mål för unionen , och en uppgift som alla parlamentsledamöter , rådet och kommissionen bör åta sig under den här mandatperioden är , såsom nämnts , att skapa området frihet , säkerhet och rättvisa .
rådet i tammerfors , motor och upphovsman till denna målsättning , föreslog vissa mål , men fem år för att utveckla avdelning iv i fördraget är för lång tid att vänta för att lösa vissa problem som brådskar .
min första tanke är att parlamentet inte bör utelämnas från de viktiga beslut som skall fattas i den här frågan och att vår delaktighet i beslutsförfarandet måste garanteras , särskilt när det gäller ett projekt för medborgarna , som kommissionären uttryckte sig så väl .
min andra tanke är att vi skyndsamt måste anta ett gemensamt system för asyl genom att godkänna gemensamma förfaranden , men framför allt genom att sätta stopp för den förvirring som nu råder mellan emigration av politiska skäl och den berättigade av ekonomiska skäl .
de sist antagna utlänningslagarna i mitt land , spanien , eller i belgien , är en larmsignal för att immigrationspolitiken skyndsamt måste införlivas .
min tredje och sista tanke rör unionens externa åtgärder när det gäller immigration och asyl .
vi varken får eller kan ge ett intryck av att unionen bara försöker skydda sig från vågen av flyktingar och ekonomiska immigranter .
vi bör välja samarbetspolitik för utveckling med våra grannar i öst och i medelhavsområdet , men detta skall göras rigoröst med ekonomiska medel och ett nära samarbete med de offentliga institutioner som samarbetar för att skydda de medborgare som får sina mest grundläggande rättigheter kränkta eller som vill emigrera för att täcka sina grundläggande behov .
avslutningsvis , när det gäller dokumentet om de grundläggande rättigheterna , så måste europas medborgare få visualisera sitt medborgarskap .
det räcker inte med euron eller sysselsättning , inte ens med säkerhet .
de behöver den &quot; europeiska själen &quot; , som en framstående spansk professor en gång sade .
herr talman ! till skillnad från vissa andra tidigare talare , vill jag ta upp uttalandena från våra portugisiska ministrar och vitorino .
orden som denna trio uttalade lät som musik i våra öron , som ceyhun sade .
som med all musik måste det vara en fin sång som är lämpligt instrumenterad .
många av oss i kammaren ser mycket optimistiskt på de kommande sex månaderna .
sången som skall spelas kommer att vara en som europas medborgare skall lyssna på , och de vill höra den rätta sången .
som beskrivits i eftermiddag kommer det ta lång tid att överrösta vissa av de obehagliga sånger som vi hört under valet till europaparlamentet och under de senaste månaderna .
amsterdamfördraget och toppmötet i tammerfors byggde på detta projekt för ett område med frihet , säkerhet och rättvisa i europeiska unionen .
ett område är emellertid oerhört viktigt och denna kammare måste delta i detta , dvs. granskning .
det finns så mycket lagstiftning - och jag välkomnar verkligen det portugisiska programmet som presenterades för oss i förra veckan - men vi måste vara helt säkra på att det granskats , att personerna i detta parlament och ledamöterna vid de nationella parlamenten och de europeiska medborgarna känner till allt i samband med programmet .
och vi måste se till att innehållet är genomförbart , lämpligt och relevant för de olika länderna .
låt mig rikta uppmärksamheten mot vissa aspekter av de resolutioner som vi skall behandla under denna eftermiddag , av vilka det hänvisats till en eller två tidigare .
jag välkomnar styrningen mot erkännandet av rättsliga system i de olika länderna och samarbetet kring brottslighet .
detta är ett område som de europeiska medborgarna med glädje kommer att acceptera .
men kommissionen och rådet måste få veta att det finns många i denna kammare som hyser betänkligheter om t.ex. eurodac-systemet .
vi accepterar rådets dominerande roll i detta sammanhang , men det finns reservationer och jag är säker på att rådet kommer att lyssna på argumentationen från de valda parlamentarikerna när de går igenom saken mer ingående .
schulz sade tidigare i dag att han inte var säker på vad en &quot; resultattavla &quot; var för något .
alla som är engelsmän eller britter eller går på cricketmatcher vet vad en resultattavla är .
en resultattavla visar resultaten - den måste vara uppdaterad , tydlig och synlig .
jag är övertygad om att kommissionär vitorino kommer att se till att detta sker .
när de sex månaderna närmar sig sitt slut , hoppas jag att musiken fortfarande spelar och att de europeiska medborgarna fortfarande lyssnar .
herr talman ! jag vill välkomna rådets ordförande och hans kollega från justitiedepartementet , costa , och tacka dem för det välkomnande de gav mitt utskott i lissabon förra veckan och de konstruktiva sammanträden vi uppskattade .
toppmötena i amsterdam och tammerfors har gett oss mycket arbete att utföra tillsammans , som det utmärkta resolutionsförslag som utarbetats av terrón visar i dag .
jag skulle vilja ta upp tre korta frågor .
den första handlar om att vi behöver ett moget samtal mellan rådet och europaparlamentet .
det är knappt sex månader sedan det genom amsterdamfördraget blev obligatoriskt för våra två organisationer att arbeta tillsammans ; vi har bedömt varandra , vi har haft några smågräl , men vi måste arbeta effektivt tillsammans .
låt oss sluta med skuggboxningen .
låt oss sluta med de omständliga charaderna och börja respektera de åtaganden som vi tagit på oss enligt fördragen och den tid det tar för en fullständigt demokratisk debatt .
låt oss delta i era diskussioner om både politik och förfaranden .
låt oss inte låtsas som om de nationella parlamenten kan utöva någon effektiv demokratisk kontroll över regeringsverksamheten inom detta område .
min andra fråga handlar om att vi behöver en kommission som har tillgång till lämpliga resurser .
vi har inrättat ett nytt generaldirektorat , ändå har detta bara 70 anställda .
det finns ett avtal om att fördubbla denna siffra , men jag har förstått att inte en enda person har anställts ännu .
vi ger kommissionen en tung uppgift , inte minst rörande utarbetandet av &quot; resultattavlan &quot; .
rådet och parlamentet måste samarbeta för att tillhandahålla de resurser som kommissionen behöver .
till sist , om debattinnehållet , välkomnar jag det faktum att ordförandeskapet placerat området för frihet , säkerhet och rättvisa högst upp på sin dagordning .
alla goda ting äro tre , i synnerhet inom vårt politikområde .
för tvåhundra år sedan var det frihet , jämlikhet och broderskap och allt gick mycket bra ända tills olika vänsterregeringar satte jämlikheten över de andra .
nu är det frihet , säkerhet och rättvisa och jag hoppas att de nuvarande vänsterregeringarna tar intryck av kommissionär vitorinos ord och motstår frestelsen att sätta säkerheten - hur viktig den är - över de precis lika viktiga behoven i samband med frihet och rättvisa .
kära kolleger ! även om det är lämpligt att erinra om de viktigaste genomförandena i den europeiska uppbyggnaden av ett område för frihet , säkerhet och rättvisa , återstår fortfarande mycket att göra .
eg-domstolens roll är fortfarande alltför begränsad och överföringen till gemenskapsnivå förblir ofullständig .
det räcker med att titta på belgiens unilaterala beslut att återupprätta gränskontrollerna .
beslutet att upprätta en stadga över de grundläggande friheterna är positivt , men det är svårt att förutse om dess innehåll och dess rättsliga omfattning , tvingande eller symbolisk , skall omfatta alla medborgare , oavsett nationalitet , eller utesluta vissa .
man kan bara beklaga den totala avsaknaden av framsteg när det gäller det europeiska medborgarskapet och politiska rättigheter för alla invånare i europa .
även om handlingsplanen från högnivågruppen syftar till att i framtiden begränsa migrationsströmmen , förbättrar dessa planer inte på något sätt situationen för de mänskliga rättigheterna , de offentliga friheterna eller den ekonomiska situationen i de berörda länderna .
vi vet att klausuler om återintagande finns i samarbets- och associeringsavtalen .
men de utgör ett allvarligt hot mot principen om icke-avvisning .
man måste också notera att dessa bestämmelser antagits inom rådet genom ett förfarande utan debatt och utan att parlamentet rådfrågats .
det grundläggande problemet är ändå ....
( talmannen avbröt talaren ) .
herr talman ! jag vill i likhet med mina kolleger välkomna rådets företrädare , såväl som kommissionsledamoten .
jag tackar dem för deras uttalanden i kammaren .
i stället för att ta upp de redan diskuterade områdena , vill jag ta upp ett specifikt ämne : narkotikafrågan och hur vi tar itu med den omfattande drogkulturen i våra samhällen .
jag vänder mig särskilt till det portugisiska ordförandeskapet och uppmanar detta att bygga vidare på en del av det fantastiska arbete som utfördes av det finländska ordförandeskapet när det gällde att utarbeta samordnade planer och åtgärder mellan medlemsstaterna .
på den internationella sidan har vi redan börjat tillämpa planer för att bekämpa narkotikasmuggling , penningtvätt osv. men vi måste föra ned det på ett mer mänskligt plan : att ge hjälp till de som försöker sluta med droger och ge dem lämpliga kontroller och lämpliga mekanismer för rehabilitering ; för det andra , att vidta samordnande åtgärder inom polisen och det rättsliga området vad gäller gemensamma straff och gemensam lagstiftning ; för det tredje , att genomföra en informations- och medvetandehöjande kampanj för yngre personer ; och en gång för alla stoppa användningen av de mycket farliga orden &quot; normalisering &quot; och &quot; skademinskning &quot; , och visa att all avmattning rörande vår beslutsamhet att se till att narkotika inte blir lagligt måste vara för medborgarnas bästa .
herr talman ! jag skulle vilja använda de futtiga sekunder talartid jag fått till att påpeka för kommissionens företrädare eller påminna honom om att regeringen i medlemsstaten belgien just nu för en politik som innebär att tusentals och måhända tiotusentals illegala invandrare blir legaliserade , kommer att få permanent uppehållstillstånd , rätt till familjeåterförening , och så vidare .
det är en åtgärd av den belgiska regeringen som är en flagrant överträdelse av schengenavtalet .
den 23 december lämnade jag in ett skriftligt klagomål om det till kommissionär vitorino .
jag skulle vilja be honom överväga det klagomålet och inom överskådlig tid tala om för mig vilka åtgärder kommissionen skall vidta för att straffa den belgiska statens överträdelse av schengenavtalet enligt artikel 226 i avtalet .
herr talman , herrar ministrar , herr kommissionär ! 1999 års skörd av beslut var verkligen riklig . så riklig , skulle jag vilja säga , att det blir svårt att ta hand om den , det vill säga att genomföra besluten .
jag syftar särskilt på rådet och på medlemsstaternas slapphet att genomföra det som man bestämmer gemensamt .
året som gick kännetecknades emellertid av flera positiva och avgörande beslut , till exempel trädde amsterdamfördraget i kraft , schengenavtalet införlivades i gemenskapspelaren , rådet beslutade i köln att utarbeta en europeisk stadga för grundläggande rättigheter och vid det extra rådstoppmötet i tammerfors förband sig medlemsstaterna att följa vissa gemensamma riktlinjer , prioriteringar och mål , med avsikten att skapa ett gemensamt område för frihet , säkerhet och rättvisa .
samtidigt som vi erkänner de framsteg som har gjorts , betonar vi , som europeiskt parlament , den ovilja som har observerats hos rådet att genomföra besluten på många områden , bristen på samsyn och , framför allt , bristen på öppenhet och samarbete med europaparlamentet .
som jag sade märker ni kanske att europaparlamentet inte är berett att spela endast observatörens roll .
det kommer inte heller att upphöra med att ställa besvärliga frågor , som till exempel om hur långt ni är beredda att gå och vilka lagstiftningsåtgärder och andra åtgärder ni kommer att vidta för att bekämpa skammen med prostitution , barnpornografi på internet , narkotikan och den organiserade brottsligheten .
kommer ni att arbeta för en gemensam asyl- och invandringspolitik ?
vad kommer ni att göra för att integrera invandrarna socialt , återförena familjer och ge tillgång till rättigheter och skyldigheter som är likvärdiga dem som gäller för medborgarna i unionen ?
kanske kommer ni att bli tvungna att överge era traditionella konservativa åsikter om flyktingar och invandrare , inför den nya demografiska ordningen som beskrivs av fn : s sakkunniga .
jag har stora förväntningar på det portugisiska ordförandeskapet .
herr talman ! jag välkomnar mycket , faktiskt det mesta , av vad som sagts under denna debatt .
men jag vill att vi iakttar försiktighet .
vi riskerar att få för många , inte för få , rättighetsstadgor i denna gemenskap : konventioner på nationell , unions- och europeisk nivå ; det är inte får få domstolar som har det sista ordet om våra rättigheter , utan möjligen för många - vi har domstolen på andra sidan floden och domstolen i luxemburg .
det finns också domstolar i karlsruhe , lissabon , dublin och edinburgh .
vi måste se till att det vi gör är förnuftigt .
vi får inte skapa förvirring och konflikter när det gäller domsrätten i samband med rättigheter , för detta skulle vara skadligt för friheten , rättvisan och säkerheten .
vi måste , kort sagt , ha och behålla högsta möjliga gemensamma standarder och hitta sätt att säkerställa dessa .
men vi måste alltid ta hänsyn till subsidiaritetsprincipen .
precis som alla andra i denna kammare vill jag ha frihet , säkerhet rättvisa .
jag vill inte se att dessa värden degenererar och skapar övercentralisering , kaos och förvirring .
fru talman , kära ledamöter !
mycket snabbt skulle jag vilja säga följande : i ledamöternas inlägg har flera frågor ställts om det portugisiska ordförandeskapet .
parlamentets talman fick oss att känna att den tid vi förfogar över är mycket kort och därför föreslår vi , jag och min kollega från justitiedepartementet , att vi objektivt besvarar alla frågor som ställs här , under mötet med det parlamentariska utskottet där vi kommer att närvara nästa vecka .
herr talman ! jag tackar rådet för såväl det muntliga som det skriftlig svaret .
effektiviteten är verkligen anmärkningsvärd .
det ger mig några sekunder extra för jag ville föreslå rådet att vi fortsätter att debattera frågan nästa gång utskottet för medborgerliga fri- och rättigheter och inrikesfrågor träffas .
då får vi tillfälle att kommentera de här svaren och uttala vår oro även inför kommissionen .
personligen är jag glad för en del av svaren , som exempelvis de känsliga frågorna om schengen eller europolkonventionen , som vi hoppas kommer att revideras , och jag gläds över justitieministerns ord i den meningen att den skall försöka underställas den dömande maktens jurisdiktion .
jag hoppas att man gör detsamma när det gäller den parlamentariska kontrollen
ärade företrädare från rådet , inom en månad kommer vi att lägga fram en resolution här i kammaren för votering .
med det goda humör som ni har visat prov på i dag , så är jag säker på att det första som kommer att hända i det här nya klimatet av samförstånd är att ni kommer att beakta resolutionsförslaget .
nästa punkt på föredragningslistan är frågor till rådet ( b5-0003 / 2000 ) .
fråga nr 1 från ( h-0780 / 99 ) :
angående : kärnkraftverk byggs på jordbävningsutsatta områden i turkiet i turkiet inträffade nyligen två jordskalv med en styrka på mer än magnitud 7 på richterskalan . det är mycket oroande att turkiet envetet tänker bygga några synnerligen kostsamma kärnkraftverk inom området akkuyu samtidigt som energin från atatürkdammarna exporteras till tredje land och eu ger ut pengar på att reparera de skador som uppstått vid jordbävningarna , i en situation där gemenskapen skär ner sin budget .
de turkiska kärnkraftsplanerna tar ingen hänsyn till de faror som kan uppstå för invånarna och ekosystemen i turkiet och omgivande länder och de inger också misstankar om att turkiets militära och politiska ledning på förhand utarbetat hemliga planer om att skaffa en teknik som skall bereda möjligheter till kärnvapenutveckling . det bör erinras att turkiet söker bygga reaktorer som är av kanadensiskt ursprung och motsvarar de reaktorer som indien och pakistan anskaffat .
vad tänker rådet göra för att kärnkatastrofer skall kunna undvikas och kärnvapenspridning förhindras till ett land som vill bli medlem av eu och som ger ut stora summor på kärnkraftsprogram men samtidigt tar emot ekonomiskt bistånd från eu ?
herr talman ! rådet vill klargöra att turkiet har skrivit under konventionen om kärnsäkerhet , vars mål ligger i linje med den oro som uttrycktes av ledamoten .
denna konvention , som trädde i kraft den 24 oktober 1996 , har just som syfte att uppnå en hög internationell kärnsäkerhet genom nationella åtgärder och genom internationellt samarbete , liksom att vid kärnkraftsanläggningarna etablera och upprätthålla ett skydd mot potentiella radiologiska risker för att skydda människor , samhälle och miljö mot skadlig joniserande strålning från denna typ av anläggningar .
konventionen omfattar som bekant också skydd mot olyckor med radiologiska konsekvenser och ett minskande av dessa effekter när den här typen av olyckor inträffar .
jag skulle dessutom vilja påpeka för ledamoten att turkiet , som ansökarland till europeiska unionen , förr eller senare , och detta är ett villkor innan anslutning - och jag tror att denna punkten är viktig - , i sin egen föranslutningsstrategi måste anta en politik som gör att landet i tid kan godta gemenskapslagstiftningen i helhet , inklusive alla bestämmelser som gäller för kärnsäkerhet .
jag skulle dock vilja tillägga följande .
med denna enhet kommer turkiet att öka sin energipotential med bara 2 procent .
det sägs emellertid att turkiet vill skaffa reaktorer av candutyp , likadana som pakistan och indien har och med vars hjälp de har framställt kärnvapen .
mot den bakgrunden måste saken undersökas , eftersom den känsliga situationen i kaukasus kan leda in många i konstiga tankebanor .
för det andra , angående anläggningarnas säkerhet .
i regioner med stor jordbävningsfara räcker det inte med att vi har starka , jordbävningssäkra hus , för vid denna slags situationer - och jag säger er detta som ingenjör - använder vi modeller för att undersöka följderna av olika faror .
vi kan emellertid inte göra modeller av kärnkraftsanläggningar i drift . det går inte .
därför kan man a priori och på förhand säga att det inte går att ha kärnkraftsanläggningar i regioner med stor jordbävningsfara .
av den anledningen , och eftersom turkiet nu står på tröskeln till europeiska unionen , måste vi hjälpa landet att bli ett säkerhetens , fredens och samarbetets land i regionen .
det är vår roll , och det är målet med min fråga .
- ( pt ) herr talman ! jag medger att de argument ledamoten framför är befogade .
det handlar i verkligheten om en mycket känslig fråga .
det är alltså en fråga , som ni förstår , som inte bara gäller turkiet i sin närhet till den nuvarande europeiska unionen , det gäller också andra stater som vi har förbindelser med genom vårt eget grannskap .
vi förstår er oro och vi kommer att ta hänsyn till den , främst inom ramen för de framtida kontakterna med turkiet när vi fastställer själva dagordningen för anslutningsstrategin för turkiet .
denna fråga hör till våra huvudangelägenheter och europeiska kommissionen kommer med all säkerhet att beakta den .
tack , herr talman och tack , herr rådsordförande !
jag är säker på att rådsordföranden är en mycket trevlig man och att han är mycket vänlig mot sin fru , sina barn och sin hund .
ni måste emellertid förlåta mig om jag är litet skeptisk rörande det svar ni just gett mig .
jag tror inte att de uttalanden som görs i rådet och omröstningsresultaten omedelbart finns tillgängliga för allmänheten .
kan ni därför , före nästa sammanträdesperiod i februari , skriva till mig och berätta var jag kan hitta denna information på allmänhetens vägnar så snart som rådet har antagit lagstiftning , i stället för att vänta på att den skall offentliggöras veckor senare som pressmeddelande .
kan ni skicka nämnda information till mig före nästa sammanträdesperiod ?
- ( pt ) herr ledamot ! jag vill först säga att jag undanber mig personliga kommentarer av det slag som ni inledde er andra fråga med och om ni kan bespara oss dessa i framtiden skulle jag vara tacksam .
i det ni framförde ger ni oss idén att kritiken mot rådet , förutom att den är formulerad på ett mycket speciellt sätt vilket vi också noterar , inte handlar så mycket om ogenomskinligheten , om vi kallar den så , i lagstiftningsprocessen , utan snarare om en överdriven öppenhet .
men jag skulle vilja säga , herr ledamot , att vi anser att resultaten av denna typ av arbete för öppenhet är klara och tydliga .
vi tvekar inte , herr ledamot , att upprepa denna information skriftligt , men vi kan inte gå längre än vad vi säger eftersom det vi säger är precis det fördraget kräver .
vi anser alltså att alla de element som rådets generalsekretariat förser allmänheten med är de viktiga element som krävs för att rådet skall fungera som lagstiftande myndighet .
jag anser att rådet inte försökte svara på min fråga .
jag frågade inte vad rådet ansåg om det förslag som kommissionen ännu inte har lagt fram , utan min fråga gäller den principiella tolkningen av artikel 255 i amsterdamfördraget .
medger den att man lagstiftar också om nationell öppenhetslag , inte bara om de tre institutioner i europeiska unionen som anges där ?
jag skulle gärna vilja ha ett svar på denna fråga .
anser rådet att man på grundval av artikel 255 i fördraget kan reglera nationell öppenhetslagstiftning , dvs. inte den som avser eu : s institutioner ?
- ( pt ) herr talman ! det svar ni fick var det svar som var möjligt att ge .
jag vill emellertid säga följande : tolkningen av artikel 255 i fördraget är en tolkning som också måste vara knuten till subsidiaritetsprincipen .
det finns för närvarande inget konkret förslag som gör det möjligt att arbeta med förordningen för denna artikel , och utan detta förslag är det inte möjligt att göra framsteg i frågan .
hur som helst , den första tolkning vi gör är att artikel 255 inte gör det möjligt att arbeta på ett sätt som påverkar subsidiaritetsprincipen .
jag är absorberad av det sätt på vilket rådet kämpar för de principer som finns i amsterdamfördraget , och som handlar om att se till att medborgarna får en bättre möjlighet att delta i beslutsprocessen .
hur gör man det när man samtidigt enligt kommissionens uttalande - det har läckt ut , så det är allmänt känt - säger att de anställdas tankefrihet sätts framför öppenheten , så att man inte kan få tillgång till arbetsdokument , rapporter , förslag osv. ?
anser inte rådets företrädare att detta försvårar ett deltagande i den demokratiska beslutsprocessen ?
fru ledamot ! den fråga ni har ställt är av största vikt och vi diskuterade den länge under senaste regeringskonferensen .
och jag vill säga er en sak : gemenskapsinstitutionernas öppenhet fungerar inte bara &quot; utåt &quot; , de fungerar också &quot; mellan &quot; gemenskapens institutioner .
det vill säga , det finns saker i formen och arbetsprocessen i gemenskapsinstitutionerna som inte är tillgängliga för andra institutioner , och det gäller inte bara mellan kommissionen och parlamentet , det gäller också mellan kommissionen och rådet .
detta ämne har alltså redan tagits upp och diskuterats flera gånger .
europaparlamentet kommer att ha möjlighet att medverka i den grupp som förbereder nästa regeringskonferens .
det är en öppen fråga .
utformningen av och den reella öppenheten i de europeiska institutionernas verksamhet är en fråga av största betydelse och det är en fråga som , enligt min mening måste analyseras än en gång , främst inom ramen för nästa regeringskonferens , detta är vi helt på det klara med , och vi menar att de ledamöter som deltar i denna förberedande grupp , får ännu ett tillfälle att ta upp denna fråga .
jag tycker att kommissionens förslag bör innehålla element för att skapa en större öppenhet i förhållande till verksamheten i de olika institutionerna , men jag menar att det alltid finns utrymme för förbättringar i denna fråga .
för vår del är vi beredda att behandla de förslag som läggs fram på detta område .
det är en väldigt viktig fråga som jonas sjöstedt och andra har ställt .
vi har en offentlighetsprincip i sverige som stärker demokratin och som ser till att det blir en bra dialog mellan medborgare , beslutsfattare och myndigheter .
vi är väldigt måna om att även eu skall gå åt detta håll , och det står även i amsterdamfördraget .
parlamentet antog ett betänkande av lööw för ett eller ett par år sedan som är väldigt viktigt i detta sammanhang .
däri varnades det för att den kommande processen skulle leda till inskränkningar i medlemsländernas offentlighet .
nu kan vi se att det kanske finns ett visst fog för denna varning från parlamentet .
jag vill fråga rådet om rådet har förståelse för denna varning , med tanke på det som vi nu har sett i arbetsdokumenten från kommissionen .
jag lyssnade med stor uppmärksamhet till det som seixas da costa sade om öppenheten och regeringskonferensen .
min fråga är om jag av det som seixas da costa sade , de intressanta sakerna om öppenheten och regeringskonferensen , kan dra slutsatsen att det portugisiska ordförandeskapet förbinder sig att arbeta och kämpa för en utvidgning av regeringskonferensens dagordning .
för undersökningen av frågan om &quot; öppenhet &quot; med avseende på institutionernas funktion kan hur som helst inte gömmas undan på något ställe och i några frågor eller i några korridorer - även om också jag inser korridorernas betydelse .
den kräver en särskilt punkt på regeringskonferensens dagordning , vilket innebär en utvidgning av denna .
- ( pt ) herr talman ! frågan om öppenhet är en fråga som naturligtvis har att göra med institutionerna .
denna regeringskonferens sätter i gång med en inriktning , åtminstone inledningsvis , på att få institutionerna att fungera bättre , särskilt med hänsyn till den önskan vi alla har om att de skall bli just mer demokratiska , öppna och effektiva .
allt detta befinner sig dock inom en allmän ram , den allmänna ramen om en gemensam acceptans av alla lösningar vi kan finna för att genomföra dessa tre önskningar .
det är uppenbart att denna öppenhet ständigt kommer att finnas med på den europeiska dagordningen och den kommer givetvis att vara med på denna regeringskonferens .
det är en fråga som det portugisiska ordförandeskapet , det kan jag försäkra er , kommer att tas upp med medlemsstaterna och företrädarna för den grupp som förbereder konferensen .
ordförandeskap bör i detta få stöd av europaparlamentets ledamöter , vilka säkerligen är beredda att stödja detta förslag .
därefter får vi se vilket resultat vi kan uppnå på ministernivå .
vi bör dock tänka på att vi just har avslutat ett amsterdamfördrag som godkändes i maj förra året , och att det där finns en mängd åtgärder för öppenhet som skall genomföras och som är på gång , och frågan är om det är för tidigt att sätta i gång ett nytt arbete om öppenhet .
jag tycker trots allt att detta är en fråga som alltid bör vara med på dagordningen , eftersom det finns en viss märkbar sensibilitet hos allmänheten angående detta , och för att det i verkligheten handlar om behovet att göra de europeiska institutionernas organ ansvariga inför medborgarna .
för vår del kommer den att finnas med .
vi får se om vi uppnår enhällighet för detta .
fråga nr 5 från ( h-0785 / 99 )
angående : förslag till förordning som anger total tillåten fångstmängd för vissa fiskarter ( i detta fall ansjovis ) för år 2000 enligt de senaste rapporterna från internationella havsforskningsrådet ( ices ) är den aktuella situationen i ices-zon viii kritisk för ansjovisbestånden .
har rådet ( fiske ) och kommissionen undersökt hur ansjovisbestånden i zon viii har påverkats av att ices-zonerna ix och x och cecaf : s ( fiskerikommittén för östra centralatlanten ) zon 34.1.1 överlåtits från portugal till frankrike ( fiskekvoterna överskrids med 5 000 ton / år ) ? har man undersökt frankrikes ansvar för den nuvarande situationen och för möjliga framtida ekonomiska och sociala konsekvenser för fiskesektorn ?
anser rådet att det är godtagbart att tillåta fortsatt överfiske som strider mot den ursprungligen fastställda totalt tillåtna fångstmängden på 33 000 ton / år , när det råder en så kritisk situation för ansjovisbestånden ?
när tänker rådet vidta några åtgärder , och vilka kommer dessa att vara , för att behandla det kritiska läge som råder för ansjovisbestånden och sätta det i samband med överlåtandet av de portugisiska kvoterna och med principen om relativ stabilitet ?
herr talman ! det portugisiska ordförandeskapet har allt intresse av att besvara denna fråga på ett fullständigt sätt , eftersom det också handlar om ett problem som berör portugal på ett positivt sätt , och jag skall förklara hur .
rådet är medvetet om den kritiska situationen för ansjovisbestånden i havet utanför kantabrien som ledamoten tar upp .
ändå ansåg de medlemsstater som utför detta fiske , det vill säga frankrike , spanien och portugal , vid det senaste rådsmötet ( fiske ) förra året , den 16 och 17 december , att tillämpningen av försiktighetsprincipen som fastställer en minskad tillåten totalfångst från 5 000 ton till 2 000 på förslag av kommissionen , var överdrivet försiktig .
man kom då fram till en kompromisslösning för att nå en balans mellan behovet att minska de biologiska riskerna , alltså påverkan på fiskbestånden , och de socioekonomiska svårigheterna som orsakas av ett begränsat fiske , med en fastställd tillåten totalfångst på en mellannivå om 16 000 ton i stället för 33 000 som var förutsett för 1999 .
en revidering planerades också i ljuset av ny information av vetenskaplig karaktär angående bevarande av arterna som man hoppas skall bli klar under första halvåret i år .
för det södra ansjovisbeståndet , i ices-zonen ix , fastställdes den tillåtna totalfångsten till 10 000 ton för år 2000 mot 13 000 ton för 1999 .
förändringarna av fiskemöjligheter mellan portugal och frankrike minskades proportionellt från 5 008 ton för 1999 till 3 000 ton år 2000 , i de franska fiskevattnen .
jag skulle vilja nämna att denna överföring inte kommer att öka fisketrycket på ansjovisbeståndet i sin helhet , inom hela gemenskapens fiskeområde .
och i enlighet med principen om relativ stabilitet , tilldelades spanien 90 procent av beståndet och frankrike bara 10 procent av fördelningsnyckeln för ansjovisfisket i havet utanför kantabrien .
utan en överföring till de portugisiska fiskevattnen , skulle den tillåtna totalfångsten i havet utanför kantabrien behöva ökas tio gånger för att ge frankrike ett adekvat fiske .
detta är skälet till att jag anser att det finns ett positivt element i portugals fall .
det är uppenbart att denna lösning skulle skada fiskbeståndet ännu mer än den risk ledamoten talade om , men vi förstår det .
herr rådsordförande ! jag måste säga att ert uttalande ingalunda har lämnat mig tillfreds .
jag förstår att portugal berörs av detta .
det är enligt min mening som ett attentat mot det sunda förnuftet och intelligensen att 80 procent av den ansjovis som fiskades i portugisiskt vatten efter avtalet mellan medlemslandet portugal och frankrike i stället börjar fiskas i biscayagolfen och att ministerrådet vidhåller att detta varken påverkar ansjovisbeståndet där eller i biscayabukten .
allt sedan 1995 har vi visat att den här omflyttningen är rena galenskapen och om portugal och frankrike vill träffa en överenskommelse så får de väl det , men ansjovisen skall fångas i portugisiskt vatten och inte i biscayagolfen .
i dag visar vetenskapliga studier att ansjovisbestånden i biscayagolfen är utrotningshotade . och nu kommer inskränkningar i de ansjoviskvoter som skall gälla för biscayagolfen .
ärade rådsministrar , jag vet inte om ni är medvetna om att ni har ett ansvar för det som hänt under de här åren men också för år 2000 när det gäller de tusentals familjer på norra delen av iberiska halvön som lever av ansjovisfiske .
- ( pt ) jag skulle vilja säga , herr ledamot , att eg-domstolen i sin dom den 5 oktober 1999 , beslutade att denna överföring , en överföring som godkändes , var i överensstämmelse med de principer som fastslås i rådets förordning 37 / 60 / 92 och främst artikel 9.1 vilken säger att medlemsstaterna kan byta hela eller delar av sina tilldelade fiskerättigheter .
domstolen uttalade också att principen om relativ stabilitet inte hade kränkts eftersom ansjoviskvoten som tilldelats spanien i underkategori 8 behölls på 90 procent och frankrikes kvot på 10 procent .
dessutom , herr ledamot , är domstolen av den åsikten att överföringen mellan portugal och frankrike inte kränker principen om rationellt och ansvarsfullt fiske i hav och levande vattendrag eftersom fisketrycket i underkategori 8 och 9 inte ökar eller innebär någon negativ påverkan för den allmänna kvoten av de resurser som tilldelats spanien .
i enlighet med detta , herr ledamot , upprepar rådet sin åsikt att utan denna överföring , skulle en hänsyn till frankrikes fiskemöjligheter göra att ansjovisfisket i biscayabukten öka .
rådet upprepar alltså , herr ledamot , sin åsikt om att fisketrycket skulle vara större och mer skadligt för fiskbestånden än den lösning som nu har valts .
konkret utgör 3 000 ton 57,5 procent av portugals fiskemöjligheter under 2000 , mot 5 008 ton , eller 73,9 procent 1999 .
dessa siffror utgör , enligt vår åsikt och rådets perspektiv , en verklig förbättring vad gäller bevarande jämfört med en nivå på 80 procent som fastställdes i rådets förordning 685 / 95 .
fråga nr 6 från ( h-0788 / 99 ) :
angående : åtgärder mot den fortgående etniska rensningen av kosovos serber och romer natos försvarsministermöte sände den 2 december 1999 ut en kraftfull appell genom vilken man kräver ett slut på den etniska rensningen av kosovos minoriteter .
europaparlamentet fördömer också i en av sina resolutioner , med hänvisning till de fruktansvärda våldshandlingar som riktats mot serber och romer , det fortsatta våldet mot den serbiska befolkningen och uppmanar de albanska ledarna i kosovo att till fullo respektera fn : s beslut nr 1244 .
i denna resolution betonar parlamentet att de tidigare förföljelserna av albaner inte kan accepteras som ursäkt för &quot; fortsatt dödande , kidnappningar , interneringar , maktmissbruk , trakasserier , hotelser , mordbränder , plundring , förstörelse av egendom och husövertaganden &quot; etc. ämnar rådet - mot bakgrund av ovanstående b ta upp frågan om finansieringen av återuppbyggnadsarbetena i kosovo till ny granskning , i enlighet med europaparlamentets krav ?
vilka övriga konkreta åtgärder ämnar rådet vidta för att få ett slut på den etniska rensningen ?
herr ledamot ! jag skulle vilja säga att jag har mycket sympati för den oro som ligger bakom er fråga .
vi delar verkligen den oro ledamoten hyser inför den hotfulla situation som råder i kosovo för de etniska minoriteterna , både den serbiska befolkningen och romerna , och som handlar om fortsatt diskriminering , förföljelser och hot på detta territorium .
rådet betonar alltid att det är nödvändigt att döma de som har begått och de som fortsätter att begå sådana handlingar rådet upprepade också , i sina slutsatser från december , att det var nödvändigt med en fullständig tillämpning av säkerhetsrådets resolution 12 / 99 och har systematiskt stött bernard kouchners arbete för att införa åtgärder som kan garantera ett effektivt skydd för minoriteterna i området , och särskilt en effektiv tillämpning av åtgärder som gör det möjligt att bevara det multietniska samhället i området .
i de kontakter vi har haft med de mest framstående politiska företrädarna för kosovos albaner , och dessa kontakter togs alldeles nyligen av den portugisiske premiärministern , har vi framhållit att förföljelserna av den serbiska befolkningen , den zigenska befolkningen och andra etniska grupper är fullkomligt oacceptabel .
detta kommer inte att tolereras och det bör genast upphöra .
detta meddelades tydligt och upprepade gånger till kosovos ledares att det internationella stödet till stor del är avhängigt av behandlingen av de icke-albanska etniska minoriteterna .
jag anser att denna punkt är av största vikt , denna känsla av förutsättning som ligger i europeiska unionens ståndpunkt kommer att vidmakthållas av rådet .
vi har stött fn-uppdragets och den internationella säkerhetsstyrkans arbete i kosovo för att förhindra nya våldsuttryck mot minoriteterna och att skydda de hotade befolkningsgrupperna .
kafor och polisen minuc ser som en av sina viktigaste uppgifter att på alla sätt få bort kränkningarna på grund av etniskt ursprung .
i detta sammanhang gläds rådet i sina slutsatser från december , åt det substantiella bidrag som europeiska kommissionen har meddelat att den skall ge indirekt till normaliseringen av situationen tillsammans med liknande bidrag från medlemsstaterna .
emellertid , herr ledamot , är rådet också medvetet om att alla medel som ges till internationellt ansvariga strukturer i kosovo inte motsvarar de som vore önskvärda , när det gäller mobilisering i de olika medlemsstaterna , och detta begränsar den effektiva handlingsförmågan när det gäller dessa strukturer .
vi kommer emellertid att koncentrera all vår uppmärksamhet på detta problem eftersom all trovärdighet för de albanska myndigheterna och strukturerna i området också beror på dessa strukturers förmåga att visa att de kan vidta åtgärder som garanterar ett multietniskt samhälle i området .
min åsikt - och allas vår åsikt , tror jag - är att portugal , landets förre president , soares , och landets regering intog en förnuftig och moderat hållning under bombningarna på balkan .
och dagens politiska uttalande om denna fråga är mycket positivt . det vill jag betona och välkomna .
trots detta finns det anledning till oro , för samtidigt som det från europeiska unionens sida finns goda och uppriktiga föresatser , är resultaten mycket små .
den senaste tiden har vi tyvärr sett en utplåning av alla minoriteter - av serber , romer , turkar , kroater - i kosovo , och vi frågar oss vad som kommer att hända .
förenta nationernas och kouchners uppdrag i kosovo är ett misslyckande .
det faktum att vi efter ett fullständigt krig som startades för att förhindra etnisk rensning nu förekommer etnisk rensning från den motsatta sidan är ett misslyckande .
av den anledningen upprepar jag min fråga , om rådet har för avsikt att vidta mer konkreta praktiska åtgärder för att diskutera dessa frågor med kouchner , som har ett mycket stort ansvar för den situation som i dag råder i kosovo .
- ( pt ) herr alavanos ! jag kan inte hålla med er om det ni säger i den sista meningen om kouchners ansvar , och jag skulle vilja urskilja två mycket viktiga nivåer : den struktur som införts i kosovo är en struktur under fn : s beskydd .
det är en struktur som europeiska unionen har gett det stöd som varit möjligt och till vilket länderna i europeiska unionen har bidragit på olika sätt .
men det finns en sak vi inte kan förneka , det är att kouchners ansträngningar för en normalisering av situationen i kosovo är oerhört positiva ansträngningar .
oberoende av om ledamoten kan tycka , vilket vi också gör , att vissa av resultaten , av skäl som inte haft att göra med kouchner , av dessa ansträngningar inte har varit så effektiva som vi alla hade önskat .
här måste vi göra en sista distinktion i ansvarsfrågan för europeiska unionen och i detta fall främst mellan rådets möjliga handlingsförmåga i detta sammanhang , och det internationella samfundets ansvar , vilket har det allmänna ansvaret för situationen i kosovo .
europeiska unionens ansvar hör alltså till ett visst bestämt sammanhang .
det är internationella samfundet , nämligen fn , som skall avkrävas ansvar för genomförandet av resolution 12 / 99 och särskilt för logiken i denna resolution och förenligheten mellan resolutionen och verkligheten .
detta är frågor vi alla bör ställa oss , men det rätta forumet för dessa frågor är fn .
herr talman ! herr rådsordförande , jag välkomnar varmt era ord att ni har för avsikt att förbättra organisationen och att det handlar om att öka myndigheternas trovärdighet .
jag tror att vi då också bör fundera över hur vi på bästa sätt skall presentera det för allmänheten .
jag frågar mig därför : finns det egentligen några idéer om hur vi kan bearbeta medierna på detta område , hur vi kan ge journalister utbildning och hur vi på ett bättre sätt kan informera allmänheten om fredlig samlevnad ?
vi har försökt att ge materiellt stöd .
vi har också försökt att på militär väg åstadkomma fred .
hur ligger det till med våra strävanden att också arbeta med psykologiska omständigheter i detta krisområde och på så sätt ge bästa möjliga stöd ?
- ( pt ) herr ledamot ! som jag sade förstår jag er oro .
jag anser att det just nu och särskilt de senaste månaderna har skett en viss positiv utveckling vad gäller de medel kouchner kan förfoga över för ett effektivt arbete .
jag minns att jag hörde kouchner under ett ministermöte med europeiska rådet i denna fråga och många angelägenheter han då påtalade angående bristande medel för att lyckas övervinna vissa problem är i dag lösta , det vill säga , han har nu fått dessa medel .
vi har framför allt två viktiga frågor : för det första , en ökad polisens resurser , vilket var en viktig fråga för att skydda civilbefolkningen , och särskilt vissa befolkningar , och ökade anslag för att främst kunna behålla vissa viktiga administrativa och operativa funktioner i processen .
frågan , herr ledamot , och det är en fråga som vi alla borde ställa , och jag gjorde det nyligen på ett diplomatiskt sätt , gäller själva karaktären på säkerhetsrådets resolution 12 / 99 .
jag vet att det är en mycket känslig fråga men vi är alla rädda att ifrågasätta den inneboende logiken i denna resolution och möjligheten att genomföra den .
vi stöder helt och hållet dess fullständiga genomförande : vi måste dock granska denna resolution - och troligen måste fn : s säkerhetsråd förr eller senare göra detta - , för att kunna bedöma , så som har skett i andra internationella strategiska scenarier , om en viss typ av agerande och en viss typ av omständighet och balans - alltså de omständigheter och balanser som ledde till att resolutionen antogs - , skall bibehållas eller ej i framtiden .
vi bör , och detta sker från europeiska unionens sida , se till att kouchner får alla resurser , och ledamoten har rätt , vi måste regelbundet och öppet förklara för våra medborgare huruvida dessa resurser används på ett bra sätt eller ej .
rådet tänker givetvis under det portugisiska ordförandeskapet komma med information i denna fråga .
herr rådsordförande ! jag är helt överens med er .
problemet är inte herr kouchner , utan den rättsliga grunden han arbetar utifrån , nämligen resolution 1244 .
jag tror därför att det är unionens ansvar , dvs. ert , men också vårt , att börja arbeta för att komma förbi den provisoriska karaktären i resolution 1244 och tänka oss ett framtida scenario för hela regionen .
jag tror att det är denna brist på definition av scenariot som åstadkommer eller gynnar de översvämningar , olyckor och mord som alavanos talat om .
avser rådet att ställa frågan om kosovos definitiva status ?
och om så är fallet , avser man att göra det i en allmän omdefiniering av regionen , och genom att så långt det är möjligt undvika att öka mikrostaterna , såsom vissa har tendens att göra , och genom att på nytt ena parterna , i detta fall kosovo och albanien ?
fråga nr 8 från ( h-0796 / 99 ) :
angående : nytt interreg-initiativ enligt kommissionens meddelande om interreg , om främjande av utveckling i städer , på landsbygden och längs kusterna , bilaga 2 punkt 1 , skall man tillåta renovering och utveckling av historiska stadscentrum med hjälp av gränsöverskridande åtgärder .
däremot framgår det tydligt att bostäder inte skall omfattas .
på landsbygden finns det många bostäder som är av historiskt intresse , exempelvis små stugor , och man bör av flera skäl bibehålla landsbygdsbefolkningarna och locka folk att bo i landsbygdsområdena . håller inte rådet med om att dessa målsättningar därför skulle kunna understödjas genom att finansiera bostadsprojekt inom ramen för interreg ?
( pt ) herr talman ! rådet , och jag skulle särskilt vilja säga det portugisiska ordförandeskapet , är oerhört medvetet om betydelsen av de problem som ledamoten fokuserar i sin fråga och jag vill säga att vi hela tiden ägnar all uppmärksamhet åt den gemensamma politiken för utveckling av landsbygden .
i detta sammanhang skulle jag vilja framhäva antagandet i maj 1999 , av ett nytt system för stöd till landsbygdens utveckling , vilket utgjorde gemenskapens referensram för en hållbar utveckling av landsbygden och det var , som ni vet , ett av de projekten inom ramen för förhandlingarna om agenda 2000 och i utvecklingen av jordbruksfrågornas hantering på gemenskapsnivå .
genom europeiska utvecklings- och garantifonden för jordbruket ( eugfj ) , är denna gemenskapens stödram inriktad på stöd till att vända tendensen till utbredning av ödemark vilket ledamoten helt befogat tar upp i sin fråga .
även europeiska investeringsfonden ( eif ) , bidrar till detta arbete med att främja den ekonomiska och sociala sammanhållningen genom att rätta till de största regionala ojämlikheterna och delta i utvecklingen och omställningen av landsbygden .
det är lämpligt att tänka på att eif har bidragit på samma sätt till främjandet av en hållbar utveckling av landsbygden som att skapa hållbar sysselsättning .
det är dessa gemenskapsinstrument i sin helhet som gör det möjligt att arbeta i en politik för landsbygdsutveckling som i dag är ett utvecklingsområde och en inriktning i den gemensamma jordbrukspolitiken å ena sidan och regionalpolitiken å den andra .
vi anser att detta , inom begreppet mångsidighet som i dag är knutet till utvecklingen av den gemensamma jordbrukspolitiken , är en av de grundläggande frågorna och eugfj : s garantisektion spelar naturligtvis här en fundamental roll .
fråga nr 9 från ( h-0798 / 99 ) :
angående : jordbruk och ordförandelandet portugal kan rådet ange ordförandelandet portugals prioriteringar för den gemensamma jordbrukspolitiken för det närmaste halvåret och de åtgärder det anser vara nödvändiga för att öka konsumenternas förtroende för jordbrukssektorn och jordbruksprodukter , efter att detta förtroende har minskat på grund av den senaste tidens hälsorelaterade farhågor ?
, rådet . ( pt ) frågan som ledamoten ställer om den gemensamma jordbrukspolitiken är en fråga som berör oss nära , och det är värt att alltid ha den med i diskussionerna i denna kammare , för vi kommer troligen att ha mycket att diskutera i detta ämne i framtiden .
under det portugisiska ordförandeskapet måste vi fortsätta debattera arbetet med den gemensamma jordbrukspolitiken , genom att anta några av de gemensamma organisationerna av marknaden med hänsyn till en harmonisk utveckling av unionens landsbygdsområden och en garanti om en positiv utveckling av jordbrukarnas inkomster , med särskild uppmärksamhet på de åtgärder som kan få följder för de små familjejordbruken .
det portugisiska ordförandeskapet kommer naturligtvis också , om den nya rundan i världshandelsorganisationen inleds under dess ordförandeskap , en sak som är långt ifrån säker , att försäkra sig om att befästa närvaron av gemenskapsproduktionen på de internationella marknaderna och en bättre balans mellan gemenskapens jordbruksprodukter som exporteras , samt bevarandet av ett mångsidigt europeisk jordbruk , vilket jag redan har nämnt .
det portugisiska ordförandeskapet kommer också att lägga vikt vid en fördjupning av politiken för livsmedelssäkerhet och detta tog den portugisiske utrikesministern och rådsordföranden för europeiska unionen , upp i dag på förmiddagen .
vi anser att livsmedelssäkerhetens roll , framför allt när det gäller folkhälsan , är en mycket viktig sak som vårt ordförandeskap skall arbeta med , det utgör för övrigt en av prioriteringarna i vårt program .
vi kommer att arbeta med detta inom fyra parallella områden inom ramen för agrifin-rådet , rådet ( hälso- och sjukvård ) , rådet ( konsumentfrågor ) och rådet ( inre marknaden ) .
det portugisiska ordförandeskapet kommer i juni i år , under europeiska rådet i santa maria da feira , också att lägga fram en rapport på detta tema , framför allt i ljuset av det som kommissionen för några dagar sedan presenterade i sin vitbok .
vi tycker att det arbete vi skall göra från och med nu för att konstituera en europeisk byrå är ett viktigt arbete för att skapa trovärdighet för den inre marknaden och för att stabilisera det egna förtroendet inom denna marknad , upplösa vissa spänningar mellan medlemsstater på detta område och till och med , varför inte säga det rakt ut , att skapa en gemensam hållning från europeiska unionens sida i sina förbindelser med tredje land på områden som handlar om livsmedelssäkerhet .
detta är det arbete vi skall försöka genomföra under det portugisiska ordförandeskapet och vi hoppas i slutet kunna presentera resultatet av detta arbete .
jag är säker på att han är medveten om det mycket allvarliga hotet mot den europeiska modellen , som grundas på familjejordbruk , i huvudsak mot de jordbrukare som sysslar med nötkötts- och fårköttsproduktion och som nu förväntas sälja sin produktion till eller under produktionskostnad .
jag vill fråga vilka nya åtgärder som rådet kan vidta för att skydda deras intressen under de kommande samtalen inom världshandelsorganisationen , i synnerhet mot den stordrifts- och industriliknande produktion som sker i förenta staterna och nya zeeland där stordriftsfördelarna gör det oerhört svårt för de europeiska jordbrukarna att skapa konkurrenskraftiga familjejordbruk och där , naturligtvis , europeiska standarder för livsmedelskvalitet inte tillämpas .
- ( pt ) jag förstår ledamotens oro fullkomligt och jag inser att det finns ett behov av vissa ansträngningar och en viss samstämmighet i frågan även inom europeiska unionen .
det är också viktigt att tänka på konsekvenserna framför allt vad gäller finansiering och ersättningar till jordbrukarna .
denna fråga är dock , som ni känner till , i händerna på europeiska kommissionen och kommer att utvecklas av kommissionen .
rådets möjlighet att ingripa på detta område är begränsat .
herr talman ! låt mig också välkomna rådets ordförande till kammaren .
men jag tror inte att han svarade på min fråga som specifikt handlade om hur vi skall ta itu med hemlöshet och bostäder , och om det portugisiska ordförandeskapet kan tänka sig att på ett aktivt sätt föra ett samtal med de icke-statliga organisationer som är verksamma inom detta område .
jag uppskattar och stöder fullständigt hans uttalande om behovet av flera strategier och ett sektorsövergripande förhållningssätt och också behovet av att bekämpa de underliggande orsakerna till utslagning , som kan leda till hemlöshet och omfatta drogberoende .
min specifika fråga handlar om problemen med hemlöshet och om det nya ordförandeskapet kan ta nya initiativ för att försöka komma till rätta med en del av de svårigheter som rådsordföranden åsyftade vad gäller stöd på mellanstatlig nivå .
jag anser att detta är ett område inom vilket europa kan spela en mycket aktiv roll , även om det bara handlar om hur utbytet av erfarenheter och bästa metoder skall gå till mellan medlemsstaterna .
- ( pt ) herr ledamot ! när det gäller ordförandeskapets möjligheter att stödja de icke-statliga organisationernas arbete , särskilt när det gäller kampen för att lösa de personliga problemen för de hemlösa , vill jag säga att denna typ av initiativ är välkomna , och vi för vår del är öppna för att diskutera möjligheter att stödja dem .
vi har samarbetat med de icke-statliga organisationerna i portugal och angående några initiativ som dessa organisationer har presenterat inom ramen för det portugisiska ordförandeskapets verksamhet och som vi knyter till alla de angelägenheter som finns i vårt eget program .
vi har inget specifikt konkret initiativ i denna fråga , vi är däremot inte låsta för tanken på att initiativ från de icke-statliga organisationerna som läggs fram för oss på detta område kan beaktas under vårt ordförandeskap .
detta , vilket måste påpekas , inom ramen för det som hör till rådets verksamhetsområde .
men vi måste förstå att allt det som handlar om kommissionens initiativrätt naturligtvis måste genomföras via kommissionen .
herr rådsordförande ! ni sade oss många saker om framtiden : vad kommissionen kommer att göra , vad ordförandeskapet kommer att göra i lissabon m.m.
och ni sade oss en sak som skrämmer mig , herr rådsordförande .
ni sade att ni i lissabon kommer att diskutera en utveckling som är mer dynamisk och konkurrensinriktad .
jag blir rädd , herr rådsordförande , för det är en sådan utveckling som leder , åtminstone delvis , till social utslagning .
jag kan inte förstå hur ni , med sådana åsikter , skall kunna ge ett svar på dessa problem .
det som jag frågade och som jag frågar igen är följande : vad är det portugisiska ordförandeskapets åsikt om de krav som kommer från t.ex. nätverken som bekämpar fattigdom och social utslagning , om fördelning av arbetstillfällen och social trygghet , om genomförandet av skattepolitiken , och då särskilt med avseende på det spekulativa kapitalet , om politiken för inkomstfördelning ?
jag skulle vilja ha ett svar på frågan om det portugisiska ordförandeskapet har för avsikt att göra någonting vad beträffar dessa saker .
- ( pt ) herr ledamoten måste förstå att ett ordförandeskaps faktiska förmåga att vända på allmänna sociala eller ekonomiska tendenser under sin period är ganska begränsad .
jag tycker att står helt klart att vår förmåga också är nära sammanbunden med vårt arbetsmetod med kommissionens initiativrätt .
jag talade det extra europeiska rådet och portugals initiativ , jag talade också om framtiden för det finns ytterligare två sätt att se på frågan om social utslagning : ett av dem är de omedelbara åtgärderna som måste vidtas för att möta dess konkreta effekter , det andra är skapandet av förutsättningar för konkurrenskraft på ett internationellt plan så att vi kan förbättra det ekonomiska taket inom europeiska unionen och få positiva sidoeffekter för problemen med social utslagning .
det portugisiska ordförandeskapet har således inga universalmedel för att under sex månader lösa de frågor som vi alltid har med oss .
vi är beredda att agera utifrån kommissionens förslag inom de områden som hör till gemenskapsbefogenheterna .
vi har givetvis både möjlighet och intresse av att få i gång alla de åtgärder som läggs fram , framför allt av icke-statliga organisationer , men också i en traditionell mellanstatlig förbindelse på detta område .
men vi måste vara medvetna om , herr ledamot , att det inte är möjligt att agera på ett område av så stor betydelse , ur ekonomiskt perspektiv , bara genom åtgärder som föreslås av ett ordförandeskap under en sexmånadersperiod .
vi tycker därför att det är klart att alla de åtgärder vi har pekat på angående strategier på längre sikt , oberoende av att vi vet att en del av de hemlösa på lång sikt kan vara döda , är de som kommer att göra det möjligt att få en hållbar politik i europeiska unionen .
det är dessa strategier som vi vill försöka bidra till på bästa möjliga sätt under vårt arbete .
fråga nr 12 från ( h-0801 / 99 )
angående : portugals ordförandeskap och utvecklingspolitiken kommer rådets sittande ordförande att uttala sig om prioriteringarna för portugals ordförandeskap när det gäller utvecklingspolitiken , lomékonventionen och hanterandet av svältsituationer ?
jag vill tacka ordförandeskapet för det omfattande svaret på min fråga , och även ministern som uttalade sig i utskottet för utveckling och samarbete förra veckan i bryssel , där han presenterade ståndpunkten .
men det finns fortfarande vissa frågor som är obesvarade .
det verkar inte finnas någon betoning på kampen mot aids i programmet. aids-situationen i afrika är nu så allvarlig att det dör fler människor i aids än p.g.a. krig .
jag hoppas att ministern kommer att lägga ned en viss tid på denna specifika fråga .
det finns tillgängliga mediciner i förenta staterna , men förenta staterna tillverkar dem inte tillräckligt billigt för de drabbade i afrika .
jag vill fråga ministern vad han tänkt göra åt situationen som håller på att utveckla sig i etiopien , där det råder torka , där skörden har slagit fel och där vi om sex månader oundvikligen kommer att vara tillbaka i det läge som rådde för några år sedan i landet , med svält och tusentals människor som dog .
samtidigt är det krig mellan eritrea och etiopien och vapenindustrin i europa är inte sen att skicka vapen , efter vilka vi skickar bröd .
- ( pt ) ledamoten måste förstå att jag först och främst inte håller med om er tolkning av min kollegas inlägg under mötet med utskottet för utveckling och samarbete , det finns inget motsägelsefullt mellan dessa ståndpunkter , snarare tvärtom .
vi kan inte i ett ordförandeskapsprogram , så vitt vi inte drabbas av storhetsvansinne , göra ett uttömmande inventarium av all möjliga och imaginära situationer för alla stora frågor som dyker upp inom ramen för internationella förbindelser .
det skulle som ni förstår vara enkelt att göra det .
det räcker med att ta en ordlista över utveckling och placera dem där , ord efter ord .
vi är tillräckligt ansvarsfulla att förstå att vi bara kan ta upp de vi har förutsättningar att klara av under vårt ordförandeskap och inom vilket - och vi bör alltid vara medvetna om detta - regeringarnas kapacitet inom rådet .
vi bör inse att det finns begränsningar vad gäller förvaltningen av de nationella vägledande programmen .
ledamoten tog upp frågan om etiopien , vilken hör till de nationella orienteringsprogrammen , men det finns som ni känner till olika gemenskapsåtgärder till kampen mot aids , och i denna aspekt har ni rätt , herr ledamot , troligen agerar inte heller usa på bättre sätt .
när det gäller politiken för utvecklingsbistånd anser jag att europa inte har något att oroa sig över av det enkla skälet att vårt agerande i denna fråga kan mäta sig med usa : s .
ledamotens fråga kom in på frågan om rustningsproblemets effekter , och det är en mer långtgående politisk fråga som jag inte tycker inryms i denna fråga men som rådet naturligtvis i framtiden kommer att ta itu med , om man anser att man skall det , och lösa genom att sätta in det i sitt speciella sammanhang .
är rådet medvetet om de sociala problem som den eu : s livsmedelsexport till u-länderna som sker till priser under produktionskostnaderna ?
har ordförandestaten för avsikt att göra någonting åt den saken ?
jag tackar rådsordföranden och framför till honom min personliga välkomsthälsning till den portugisiska regeringens ordförandeskap .
tillåt mig att tala om för honom hur vältalig och kunnig han är om de europeiska frågorna .
eftersom rådet erkänner kulturens stora betydelse som ekonomisk handelsvara , borde det , enligt min åsikt , visa det även i praktiken . och jag är rädd för att ursäkten att kultursektorn styrs av subsidiaritetsprincipen , och följaktligen är de nationella regeringarnas ansvar , är ett svepskäl .
för den fråga som jag ställde och som förblev obesvarad är varför rådet , liksom för övrigt också kommissionen , när europaparlamentet begär ökade anslag för att finansiera europeiska unionens kulturprogram , regelmässigt minskar dessa och ibland till och med avslår dem helt . det visar i praktiken rådets ointresse för kulturen , trots rådets motsatta försäkringar om att det tillskriver kulturen stor betydelse .
jag skulle alltså vilja fråga rådet om det är berett att från och med nu stödja kulturen , med samma iver som det subventionerar bananerna , humlen , korna och cannabisen .
ordet går till dimitrakopoulos för en ordningsfråga .
jag vill bara informera er om följande : i morse förövades ett attentat i madrid .
en bomb hade installerats i en bil . en person har dött .
jag vill bara å min grupps vägnar än en gång fördöma dessa terroristhandlingar .
tack så mycket , fru fraga .
vi har faktiskt blivit informerade om den tragiska händelsen .
än en gång bestraffas tyvärr det spanska samhället av dessa mordiska terrorister .
ordförandeskapet noterar era ord med särskild intensitet eftersom ordförandeskapet vid dagens sammanträde också är spanskt .
jag förklarar europaparlamentets session återupptagen efter avbrottet den 21 januari 2000 .
fru talman ! tillåt mig påminna om att i morgon är det två år sedan katastrofen i cermis .
för två år sedan kapade ett amerikanskt flygplan från natobasen i aviano under en övningsflygning på låg höjd - under den tillåtna säkerhetsgränsen - linorna till en linbana i cavalese i italien och orsakade över 20 europeiska medborgares död .
alltsedan dess väntar offrens familjer , som inte har kunnat söka tröst i någon rättvisa eftersom den ansvarige piloten inte har fått något straff , på att få åtminstone ekonomisk ersättning från usa .
jag vill därför uppmana parlamentets talman och rådets ordförande att hos de amerikanska myndigheterna utverka en omedelbar ersättning i enlighet med de rättigheter som offrens familjer har .
tack , fru angelilli !
efter den begäran jag erhållit från flera politiska grupper och efter den talmanskonferens vi just haft , föreslår jag en debatt på en och en halv timme om en aktuell och brådskande fråga av större vikt , i enlighet med artikel 50 i arbetsordningen , om unionens reaktion på regeringsförhandlingarna i österrike .
om ni beslutar att föra upp denna debatt på föredragningslistan kommer den att inledas av rådets ordförande seixas da costa och kommissionens ordförande romano prodi .
vill någon uttala sig för detta förslag ?
finns det någon kollega som vill uttala sig emot detta förslag ?
fru talman ! jag vill uttala mig emot av principskäl som förefaller mig fullständigt grundläggande , eftersom det handlar om att respektera fördragen , bl.a. artikel 7 i amsterdamfördraget .
fru talman , kära kolleger ! vi har hittills trott att europeiska unionen , enligt bestämmelserna i rom- och parisfördragen genom vilka gemenskaperna grundades , och som sedan blev unionen , var en sammanslutning av fria , oberoende och suveräna stater .
även om ett stort antal förändringar gjorde att vi betvivlade detta , har vi ändå ansett att detta var fallet och nyligen hänvisade man återigen till subsidiaritetsprincipen , även om det var halvhjärtat . fru talman !
det förefaller emellertid i dag uppenbart att om man inleder den debatt som ni och talmanskonferensen ber oss att inleda , på grundval av artikel 50 , skjuter man en fruktansvärd bräsch i principen om frihet , staternas suveränitet och regeringarnas fria sammansättning , som är resultatet av demokratiska val , och då kan i morgon en annan majoritet i parlamentet lägga sig i bildandet av en regering som ändå är resultatet av fria , regelrätta , fredliga och demokratiska val inom en medlemsstat .
om ni ratificerar ...
herr gollnisch ! ursäkta mig , men ni har bara en minut .
jag vet att ni alltid är noga med att arbetsordningen skall respekteras .
fru talman ! jag trodde att jag hade tre minuter .
om ni ratificerar denna utveckling ratificerar ni utvecklingen av en union i riktning mot en organisation som kommer att bryta mot suveräniteten och friheten för medlemsstaternas nationer , och vi har då inget annat val än att utträda ur en sådan union .
regeringsförhandlingar i österrike
nästa punkt på föredragningslistan är debatten om regeringsförhandlingarna i österrike .
jag ger genast ordet till rådets ordförande .
fru talman ! min grupp välkomnar denna debatt för den är betydelsefull .
detta är första gången i det moderna europeiska projektets historia som vi börjar se ett parti från extremhögern integreras i politiken .
det är djupt oroande .
fpö hävdar att om man läser deras litteratur och deras programförklaring finns där mycket som man skulle kunna känna sig delaktig i .
så är det kanske men låt mig i dag föra till protokollet den långa och svåra upplevelse som vi liberaldemokrater genomgick med österrikiska fpö inom vår familj liberal international .
så tidigt som 1986 hade vi anledning tro att jörg haider inte var en man vars principer eller inställning överensstämde med anständighet och modern liberalism .
i november 1991 efter en lång intern debatt inom liberal international och många besök i wien för att diskutera frågor avstängde vi temporärt fpö som medlem och i juli 1993 uteslöt vi dem .
( applåder ) vi uteslöt dem då och vi fortsätter att förkasta det som haider står för nu .
låt mig berätta för er vad vi lärde oss under denna långa erfarenhet .
det fanns många bland oss som sade &quot; läs texten &quot; .
det fanns många fler bland oss som sade &quot; läs undermeningen &quot; , &quot; se på kontexten &quot; .
ord som används i politiska sammanhang kan vara uppviglande , kan vara upphetsande eller försonande .
vi ansåg att jörg haider , som ordvrängare , har varit en röst för rasism och för främlingsfientlighet .
han är en man som spelar på rädsla och som har utnyttjat människors sårbarhet .
det är därför denna debatt är viktig - att markera att när man integrerar extremism händer något mycket omvälvande i europa i dag .
jag skyndar mig att tillägga att vårt gräl inte gäller det österrikiska folket .
vi respekterar det österrikiska folkets rätt till sin egen demokratiska process .
vi försvarar det österrikiska folkets rättigheter och konstitutionella privilegier , men vi här i europaparlamentet har en skyldighet att påminna oss om våra grundläggande principer enligt artikel 6 i fördraget - principerna om frihet , demokrati och respekt för mänskliga rättigheter .
varje rättänkande person i denna kammare anser att dessa är universella och odelbara principer utan hänsyn till färg , klass eller tro .
vi måste värna om och försvara dessa rättigheter och samtidigt tala om för det österrikiska folket : vårt gräl gäller inte er .
beträffande det portugisiska ordförandeskapets initiativ vill jag framföra att vi stöder andemeningen och det politiska syftet bakom det .
det är kanske inte ett perfekt initiativ i dess utformning men vi inser , herr ordförande , att dess grund är idealism och av det skälet är vi benägna att stödja det .
jag delar ordförande prodis uppfattning att gemenskapens metod är att föredra och vi måste titta på artiklarna 6 och 7 i fördraget .
i artikel 7 nämns möjligheten till tillfällig uteslutning i händelse av allvarliga och återkommande brott mot våra grundläggande principer .
vi måste som institutioner hitta ett sätt att tillämpa och visa vad detta betyder , så att det får en verklig mening och innebörd .
därefter kan vi arbeta tillsammans i enlighet med gemenskapens metod för att driva ut denna cancerböld mitt ibland oss .
fru talman , jag vill säga några ord till schüssel .
schüssel är en man med ett hedersamt rykte i europeisk politik .
han avser nu att rida in i regeringen på ryggen av en politisk tiger .
herr schüssel , ni tar på er ett mycket tungt , personligt , nationellt och europeiskt ansvar .
det ansvaret , som ni herr schüssel nu tar på er är att respektera ordalydelsen och andan i de europeiska fördragen .
slutligen , fru talman , detta är en debatt som berör kärnan för våra demokratiska principer och institutioner och påminner oss om att priset för frihet är evig vaksamhet .
på denna kontinent , av alla platser , och mot bakgrund av vår erfarenhet av hatisk rasism som vi utstått tidigare och till så stor kostnad måste vi hävda att dagens debatt inte handlar om att hindra en stats suveräna rättigheter .
det är ett hårdnackat krav från de demokratiskt valda i denna unions institutioner att vi som européer inte kan tillåta att man vrider tillbaka klockan .
fru talman , kära kolleger ! i dag är det hyckleriet som står på dagordningen .
vi har ett råd som lyckats strunta i fördraget och använda en metod som helt ligger utanför artikel 6 och 7 och som , vid fall av allvarliga och långvariga brott , gör det möjligt att döma en stat .
i detta fall föreligger inte allvarliga och långvariga brott i österrike .
det finns risker - det är vi alla medvetna om - men det förekommer absolut för närvarande inget som helst vare sig allvarligt eller långvarigt brott .
om man skulle tillämpa kriterierna i artikel 6 och 7 , om man skulle tillämpa kriterierna från köpenhamn på våra institutioner , på europeiska unionen , skulle denna europeiska union mycket sannolikt inte kunna bli medlem , på det sätt som man kräver av länderna i central- och östeuropa .
och om vi talar om allvarliga och långvariga brott , kan vi kanske tala om vissa medlemsstater , vi kan tala om italien och frankrike , det första respektive tredje land som dömts av europarådet , av domstolen i strasbourg .
vi kan , kära belgiska kolleger , tala om belgien , om dutroux-affären , tiotals och åter tiotals barn som rövats bort , torterats , våldtagits och mördats av personer från detta land och där undersökningarna fortfarande har kört fast .
kära kolleger ! vi skulle med en tredjedel av ledamöterna kunna tvinga rådet och kommissionen att ifrågasätta detta .
vi skulle själva kunna ifrågasätta det faktum att österrikarna förkastar tio år , tretton år av &quot; partikrati &quot; som korrumperat och fått ett land - österrike - att ruttna på samma sätt som det är på väg att korrumpera och låta länder som italien , belgien och andra av unionens medlemsländer ruttna . kära kolleger !
vi skulle verkligen kunna fråga oss varför 76 procent av de belgiska medborgarna inte har något förtroende för rättvisan i sitt land , 56 procent av de franska medborgarna inte har något förtroende för rättvisan i sitt land och 53 procent av de italienska medborgarna absolut inte har något förtroende för sin rättvisa ...
( talmannen avbryter talaren . )
fru talman ! min grupp , edd , och i synnerhet mitt parti , är mycket oroade av denna debatt .
vi kan inte stödja och vi stöder inte på något sätt haiders åsikter och politik och vi beklagar hans hänvisningar till tredje riket .
men vi beklagar dock det faktum att ert parlament överväger att blanda sig i en vald regerings politik i något som helst land , särskilt ett som är en del av europeiska unionen .
mitt parti hemma är verkligen inte rasistiskt , men vi godkänner inte europeiska unionens princip eller inblandning så lätt .
kommer ni att blanda er i politiken i storbritanniens parlament om vi blir valda ?
fru talman ! österrikes folk har talat genom att välja haider till sitt parlament .
jag tror de gav honom 28 procent av rösterna , så det kommer att bli en koalitionsregering .
fru talman , får jag föreslå att ert parlament väntar och ser om haiders parti kommer att påverka det landets politik .
då och först då kan ni bedöma om mänskliga rättigheter påverkats .
ert parlament kan överväga lämpliga åtgärder för att lösa den situationen och då , fru talman , först då kan ert parlament överväga att blanda sig i konstitutionella frågor i ett av europeiska unionens länder .
fru talman , som ledamot från det österrikiska liberala partiet respekterar jag den oro som vissa kolleger känner för den demokratiska utvecklingen i österrike .
ni kanske förvånas över min reaktion när jag säger att jag förstår att man är särskilt känslig och ifrågasätter österrikes respekt för de mänskliga rättigheterna och dess ansvarskännande gentemot det egna förflutna och i fråga om den demokratiska stabiliteten i landet .
österrike måste själv ta ansvaret för den ofta tvivelaktiga image som det med rätt eller orätt har i utlandet .
våra regeringars vägran under många år att erkänna vår delaktighet i andra världskrigets fasor , och deras vägran att rättmätigt gottgöra de judiska offren och tvångsarbetarna , har väsentligt bidragit till denna negativa bild .
nu har detta fpö ( österrikiska liberala partiet ) på grund av det uppdrag de fick vid valet den 3 oktober 1999 , när den gamla regeringen valdes bort , gått in i en regeringskoalition med övp ( österrikiska folkpartiet ) .
detta är den rättighet som medborgarna i en stat har , eftersom det är grundprincipen i en demokrati .
efter att samtalen mellan spö och övp misslyckats försökte socialisterna bilda en minoritetsregering och bad fpö om deras stöd .
vi erbjöds tre ministerposter - det kan ni se i tidningarna - just detta parti som här betecknas som fascistiskt !
när vi plötsligt avvisade detta erbjudande , började en våldsam hets och propaganda , som vi hittills inte kunnat förstå .
fpö är ett parti som länge varit etablerat inom den österrikiska politiken .
det tillsätter ministerpresidenten i ett av de nio förbundsländerna och deltar i alla andra regeringar .
varför , frågar sig många österrikare i dag , tolkas deras demokratiska beslut plötsligt som ett uttryck för en fascistisk inställning , varför har hetsen börjat just när de liberala avvisade stödet från en socialdemokratisk minoritetsregering ?
här ägnar man sig åt ett fördömande som gör den hemskaste epoken i den europeiska historien till ett politiskt spektakel - utan att gå in på vårt program .
det äcklar mig , när några av våra motståndare utnyttjar miljoner människors död i koncentrationslägrens gaskammare till billig propaganda , vilket exempelvis den italienske ledamoten bertinotti gjorde , när han i går i italiensk tv anklagade haider för att förneka förintelsen .
ni borde skämmas , herr kollega !
även om alla era politiska argument tar slut , har ni inte rätt att använda de mördade personerna för er billiga propaganda .
ni förvandlas här inte till någon antifascist när ni betecknar en demokratiskt vald politiker som nazist !
tvärtom , ni hånar de verkliga offren för nationalsocialismen och bagatelliserar de fascistiska diktaturerna .
ni agerar på grund av era egna fördomar , ni avstår från all politisk diskussion och agerar just på det sätt som ni påstår att ni bekämpar .
attacken mot österrikes nya regering , försöket att påverka politiken i ett medlemsland är en förolämpning av den österrikiska befolkningen .
därför är vi tacksamma för kommissionens speciella hållning .
i de nya koalitionsavtalen handlar det om en demokratireform , oppositionens rättigheter och plikten att lämna skadestånd åt tvångsarbetarna .
fru talman ! det här är ett historiskt ögonblick eftersom det nu äntligen står helt klart för oss alla att europeiska unionen allt eftersom utvecklats till en värdegemenskap .
vi inser detta nu när en medlemsstats regering håller på att få ett parti som veterligen inte respekterar dessa värden .
jag vill också konstatera att de fjorton medlemsstaternas ställningstagande från rådets sida var berättigat , eftersom det här på sätt och vis också handlar om sammansättningen på europeiska unionens regering , vilket gör att den här frågan angår även rådet . det är inte enbart österrikes interna angelägenhet .
i egenskap av parlamentsledamöter måste vi särskilt betona att det arbete som inletts för att förstärka de grundläggande rättigheterna t.o.m. är viktigare än förut .
det är viktigare än förut att respekten för och okränkbarheten hos de mänskliga rättigheterna samt minoriteternas rättigheter , alla de människors rättigheter som bor i europeiska unionens område , är en väsentlig del av europeiska unionens rättsstatsprincip , och därför måste också stadgan för de grundläggande rättigheterna göras juridiskt bindande .
den får inte enbart förbli en förklaring .
lika viktigt är det att stödja österrikes demokratiska krafter , ingen av oss vill ju isolera österrike .
vi vet att majoriteten av österrikarna respekterar dessa värden .
de har också demonstrerat ; alla demonstrationer har inte ägt rum utanför österrike .
det är säkert också många väljare som röstat av protest , som länge velat ha en förändring i den österrikiska politiken .
enligt min mening skall parlamentet stödja dessa demokratiska krafter .
jag vädjar också till österrikes president att han än en gång skall undersöka alla de möjligheter som finns att bilda en regering bestående av demokratiska krafter .
fru talman , kära ledamöter ! jag vill bara understryka värdet av den hållning som vår gruppordförande , francis wurtz , påminde om för ett tag sedan .
jag uppskattar uttalandet från rådets ordförande och ståndpunkten från de 14 medlemsländerna som vägrar att ha officiella kontakter med den österrikiska regeringen så länge som jörg haiders parti ingår .
det faktum att vi instämmer i detta blir desto viktigare eftersom vi , som bekant , har en kraftigt avvikande uppfattning när det gäller den politik som bedrivs av europeiska unionen . detta gäller den ekonomiska och sociala politiken , det demokratiska underskottet , det faktum att unionens medlemsstater deltog i det dramatiska kriget på balkan .
detta vårt avståndstagande understryker ännu mer betydelsen av vårt instämmande i dag : det är något exceptionellt , för faran för att ett irrationellt och neonazistiskt parti återuppstår i europa är exceptionell .
den risken gäller inte bara österrike , den gäller hela europa .
vi talar om oss själva , inte om österrike .
vi känner till de sociala faktorer som samverkar med arbetslösheten och osäkerheten , till att förstärka tendenserna i den riktningen . vi känner till de kulturella orsakerna - främlingsrädsla , rasism - men vi kan inte avstå från att i oförmågan och den bristande viljan från extremhögerns sida göra upp med nazismen och peka på risken för att det uppkommer en explosiv blandning i europa .
jag talar om alperna , om alla våra länder . vi håller på att skapa förutsättningar som kan leda till att det uppkommer en fara för demokratin och det europeiska samhället .
ordförandeskapets uttalande visade att man är medveten om det dramatiska i situationen .
europa visar att man inte har glömt auschwitz . europa möter ett spöke .
men nu måste vi vara konsekventa i våra handlingar , och den första att vara konsekvent borde vara kommissionen , som i stället här har visat prov på en oklarhet och en brist på stadga som gör ordförandeskapets ståndpunkt ännu mer värdefullt .
detta är den ändring vi måste kräva i kommissionens åtgärder .
fru talman , kära kolleger ! i den grundläggande demokratiska principen om respekt för de mänskliga rättigheterna och folkens frihet och suveränitet , mot all gammal eller ny fascism , nazism eller kommunism , och med tanke på att samtliga föregående talare har talat om det österrikiska folkets suveränitet , så ser vi i dag hur denna suveränitet förnekas av just detta parlament .
när man läser det österrikiska liberala partiets partiprogram så finner man där ingenting som rättfärdigar anklagelserna om ett attentat mot principerna om frihet , demokrati och respekt för de mänskliga rättigheterna , de principer om grundläggande friheter och om rättsstaten som framhålls i artikel 6 i unionsfördraget .
låt mig i stället rikta er uppmärksamhet på det faktum att den tjänstgörande ordföranden , som var så kritisk när det gäller österrike , nyligen överlämnat invånarna i macao till den demokratiska kinesiska folkrepublikens överhöghet .
men kanske är det i dag , för att stärka demokratin inom unionen , lämpligt att isolera österrike , kriminalisera ett parti som valts på demokratisk väg av det österrikiska folket och i stället släppa in det turkiet som styrs av de grå vargarna i europa .
fru talman , ärade ledamöter ! det är en högst allvarlig fråga vi diskuterar .
det handlar om inte mindre än närvaron av en politisk makt i en medlemsstats regering , en makt vars lärosatser och principer är oförenliga med unionens föreställningar och moral som är heliga i de fördrag som unionen bygger på .
en genomläsning av artikel 1 i kapitel 4 i det österrikiska populistiska partiets program kan uppröra vilken demokrat som helst .
accepterandet av den etniska gruppen som en avgörande faktor för en nation och påståendet att en folkgrupp är överlägsen alla andra , så som det påstås där , väcker gamla spöken till liv från ett århundrade som vi just har lämnat bakom oss , och som av vissa historiker betecknas som skräckens århundrade , en skräck som till vår bestörtning åter aktualiseras av den oacceptabla filosofin i haiders politiska program .
naturligtvis är det österrikiska folket ett självstyrande folk och naturligtvis skall vi respektera principen om icke inblandning i en medlemsstats inre angelägenheter .
men det är inte det som är problemet .
problemet är huruvida unionen kan förbli likgiltig inför bildandet av en regering i en medlemsstat , där ett parti med sådana drag ingår .
vårt svar på denna avgörande fråga är nej .
( applåder ) bortom alla strategiska och taktiska överväganden , bortom alla eventuella rättfärdiganden som man gör på grund av främmande beteenden , bortom allt sådant , och oberoende av partiintressen och valtider , vill den spanska delegationen inom europeiska folkpartiets grupp i parlamentet , helt i överensstämmelse med det spanska folkpartiet och spaniens regering , uttrycka sitt stöd för uttalandet av rådets portugisiska ordförandeskap den 31 januari , vad beträffar dess innehåll , ton och konsekvenser .
konrad adenauer sade vid något tillfälle - och han visste vad han talade om - att det säkraste sättet att lugna ned ett odjur är att låta dig slukas .
historien är en provkarta på sådant som hade kunnat undvikas .
därför , fru talman och kära kolleger , måste unionen och detta parlament ge tydliga signaler om att vi avvisar detta intoleransens , främlingsfientlighetens och totalitarismens odjur , för att bara nämna några av de misstag på den långa lista över avsägande av ideal , avståenden och opportunism som markerat europas förflutna och som vi har fått betala ett högt pris för .
fru talman , kära kolleger ! vår union konstruerades kring tanken : &quot; detta får aldrig hända igen &quot; , och detta betydde &quot; aldrig mer främlingsfientlighet , läger , antisemitism , aldrig mer någon bitter nationalism eller några krig &quot; .
europeiska unionen har inget annat syfte än viljan att överträffa denna fruktansvärda historia från det tjugonde århundradet som , i hjärtat av europa , dödade hela idealet om humanism och som i dag fortfarande är högst aktuellt .
det är inte sant när man säger att när en regering bildar allians med nyfascister , någonstans i europa , är det bara ett problem med nationell suveränitet .
vår union är inte någon sammansättning av stater-nationer som gör arrangemang sinsemellan för att förbättra sitt öde .
det är en ödesgemenskap där alla demokrater tillsammans , när det viktiga ifrågasätts , när värderingar ifrågasätts , måste stå enade för att finna lösningar så att misstagen inte återupprepas .
vi måste ta lärdom av det förflutna .
under trettiotalet valdes adolf hitler demokratiskt , även om det var med minoritet , många tyckte att det inte var så farligt och , herr poettering , i mitt land ansåg ett antal män och kvinnor till höger , men kanske också på annat håll : &quot; hellre hitler än folkfronten &quot; .
de föredrog sina lokalpatriotiska trätor framför det viktiga , och katastrofen var ett faktum .
vi måste reagera snabbt , kraftigt och enat . herr poettering !
jag skulle ha velat höra er tala till den österrikiske presidenten eftersom vi vet att han i dag är mycket generad över denna smutsiga allians som ingåtts av en regering .
vi måste alltså reagera snabbt och kraftigt .
naturligtvis innehåller fördraget en spärr när handlingarna blir outhärdliga , och jag höll nästan på att säga &quot; irreparabla &quot; .
historien har lärt oss att fascisterna börjar med att ge ros och ris : först ris , i de populistiska och främlingsfientliga talen , och sedan ros för att göra sig presentabla i institutionerna och successivt infiltrera dem , fördärva dem , ända till den dag de skrider till handling .
och den dagen är det för sent .
fördraget innehåller därför spärrar ; men vi är inte där ännu ; i dag måste vi förhindra att vi kommer så långt som till dessa spärrar .
vi måste därför finna en politisk lösning .
i det stöder jag rådets förslag och jag beklagar en viss ömtålighet , en viss slapphet från kommissionen som ändå borde vara beslutsamt vaksam dag för dag , för fascisterna räknar med demokratins slapphet , de räknar med tiden för att slita ut oss och de hoppas slutligen kunna göra sig gällande .
vi måste därför reagera snabbt .
om vi i dag inte starkt stöder rådet kommer historien att döma oss och säga : de har genomfört ett politiskt münchen .
fru talman ! jag gläder mig över att den stora befolkningsmajoritetens vilja respekteras i österrike och att , ur min synpunkt , demokratin vunnit en mycket viktig seger i och med den här regeringsbildningen .
det måste stå alldeles klart : ett europa som utvecklas som en sorts &quot; big brother &quot; som på stalinistiskt sätt och med stalinistiska metoder vakar över vänsterns political correctness i den ena eller den andra medlemsstaten , ett sådant europa undanber vi oss verkligen .
den europeiska demokratin och den österrikiska demokratin behöver inte ta emot lektioner från någon annan och särskilt inte från en belgisk regering , till vilken av vapenhandlare finansierad korruption hör . en belgisk regering som utsett ordföranden för ett sådant av domstolarna korruptionsdömt parti till ledamot av europeiska kommissionen .
vi tackar i dag österrikes befolkning för den här demokratiska segern som är viktig för alla folk i europa och för var och en som förespråkar frihet och yttrandefrihet .
fru talman , rådets företrädare , herr kommissionär ! för en vecka sedan avslutades i stockholm den stora internationella förintelsekonferensen .
dess syfte var att bekämpa glömskan och det onda i dagens samhälle som uppträder i form av främlingsfientlighet och nynazism .
det vore ett hån mot idén bakom denna konferens och hela det internationella samfundet att i dessa tider inbjuda ett nazistflirtande och främlingsfientligt parti i eu : s institutioner .
för det andra vill jag säga att vi måste vara konsekventa mot oss själva och våra värderingar .
vi kräver av kandidatländerna och av samarbetsländerna i loméavtalet att de skall respektera mänskliga rättigheter och visa tolerans gentemot nästan .
vi måste göra detsamma mot oss själva .
det är därför vi reagerar mot detta smusslande som pågår i österrike .
det går inte att fortsätta som om ingenting har hänt .
vi står inför en vattendelare i unionen .
unionen är inte bara en ekonomisk gemenskap , utan det är en värdegemenskap som vi tar på allvar .
någonting har hänt : unionen håller på att få ryggrad och själ .
vi är bekymrade . vi , det är de belgiska kristdemokraterna och lyckligtvis väldigt många andra kolleger med oss .
den koalition som håller på att bildas i en av medlemsstaterna är absolut en österrikisk angelägenhet men det hela har utan tvivel även en europeisk dimension .
vad binder oss samman i europa .
i första hand värdena och principerna om frihet , demokrati och respekt för de mänskliga rättigheterna .
ordföranden för det österrikiska liberala partiet , haider , har flera gånger visat att han inte tillräckligt högt värderar ens de grundläggande formerna av diplomatisk artighet .
han är en farlig man .
de kristdemokratiska partierna i mitt land har för länge sedan valt , och håller fast vid , att visserligen lyssna till de högerextremistiska väljarnas protester men att aldrig förhandla med de högerextremistiska ledarna .
värden måste komma före makt .
därför beklagar vi det som sker i österrike .
vi är till och med skakade av det .
vi är mycket besvikna .
vi uppmanar övp att i sista hand ändå undersöka andra lösningar .
vi fortsätter att påminna om artikel 6 i fördraget .
vi fortsätter kämpa mot banaliseringen av den extrema högern .
om koalitionen ändå blir av så uppmanar vi våra kolleger i övp att både i program och i ord och handling garantera att de principer och värden som utgör grunden för den europeiska integrationen respekteras .
fru talman , mina damer och herrar , kolleger ! det vilar ett stort ansvar på österrike .
( en ) fru talman ! där jag kommer från säger man &quot; en walesare har tre tillfällen &quot; och tre gånger , vilket jag tror ni kommer att upptäcka under den debatten , framförde jag min önskan att kortfattat lämna synpunkt på vad som har varit en utmärkt och vid flera tillfällen känslig debatt .
först och främst vill jag framföra mitt tack på ordförande prodis vägnar och mina kollegors i kommissionen för det stöd och samförstånd som flera ledamöter av kammaren visade för kommissionens ståndpunkt i det uttalande som vi gjorde i går .
jag måste naturligtvis även reagera på det faktum att man under debatten gjorde anspelningar på - och jag använder några av de ord som användes - tvetydigheten , eftergivenheten och vekheten i kommissionens yttrande .
jag känner mig förpliktad att till denna kammare framföra att det finns ingen tvetydighet eller vekhet eller eftergivenhet i det yttrande som gjordes eller de åtgärder som kommissionen vidtog i denna fråga .
vi hänvisade i vårt uttalande i går morse , liksom ordföranden gjorde i eftermiddags , uttryckligen till det faktum att vi delar den oro som fjorton medlemsstater framförde i sitt uttalande i måndags .
för det andra , påpekade vi i mycket specifika termer att vi kommer att arbeta nära och tillsammans med alla medlemsstater för att granska situationen och dess utveckling i österrike .
för det tredje , vi förklarade mycket klart att vi utan rädsla opartiskt kommer att hålla fast vid principerna och bestämmelserna i artikel 6 i fördraget och att vi skall göra vad som ankommer på oss enligt artikel 7 i fördraget för att säkerställa att dessa principer för frihet och demokrati och grundläggande fri- och rättigheter upprätthålls .
det finns alls ingen eftergivenhet , vekhet eller tvetydighet i något av detta .
och när jag säger att kommissionen intog denna ståndpunkt innefattar jag min kära kollega franz fischler , som kommer från österrike och som återigen bevisade sin integritet och sin oberoende ställning som ledamot av europeiska kommissionen under ed genom att delta i det uttalande som vi gjorde i går morse .
var och en som därför bjuder in franz fischler till sitt hem för att av någon anledning förklara det faktum att han är av österrikisk nationalitet bör granska sina egna motiv i samband med en debatt som nödvändigtvis har skymts av hänvisningar till främlingsfientlighet och även mer farlig ondska i denna värld .
jag säger det i vänskap och vördnad för min vän och kollega franz fischler .
får jag också tillägga , fru talman , att förståelsen hos ordförandeskapet , det portugisiska ordförandeskapet , för vår ståndpunkt mycket klart bekräftades av da costa när han sade , och jag citerar honom , att &quot; portugal och övriga medlemsstater önskar säkerställa att gemenskapsmaskinens arbete inte störs av den nuvarande situationen &quot; .
det är förvisso i allas intresse .
för att kunna garantera att fördraget efterlevs och att vi håller vad som beskrevs som gemenskapsmaskinen i gång följer vi det tillvägagångssätt som lades fast i vårt uttalande i går .
vi skall fortsätta att göra det , fru talman , på ett opartiskt sätt .
det är vår plikt .
det är också en fråga om övertygelse .
min sista punkt är följande .
vi inser innebörden i denna viktiga debatt .
det finns flera personer här som liksom jag själv under många år tidigare blivit vana vid haiders stötande uttalande , främlingsfientligheten i många delar av hans politik och den strategi han utvecklat att omväxlande göra aggressiva uttalanden och sedan framföra ursäkter , ibland påföljande dag .
vi inser det och vi kommer även ihåg det dåliga och selektiva minne han ibland visar om nazismen .
och när vi minns det , som så många andra runt om i denna kammare , väcks naturligtvis mina och mina kollegors instinktiva känslor till liv .
men kommissionen måste agera på grundval av värderingar och lagar och inte bara på grundval av instinkter .
det är därför vi kom fram till vår slutsats i går morse .
det är därför vi håller fast vi den slutsatsen medan vi fortsätter att upprätthålla principerna och lagarna .
utan vekhet , utan eftergivenhet , utan tvetydighet men till nytta för hela unionen och varje medlemsstat i unionen och dess folk .
vi skall fortsätta att göra det energiskt och konsekvent och som cox sade i debatten , &quot; ovillkorligen med hög bevakning &quot; .
jag undrar , då da costa har lyssnat till dessa inlägg långt bak i kammaren , om herr kinnock kan bekräfta att kommissionen stöder den åsikt som da costa klart fastslog i dag och som även fastslogs i ordförandeskapets nyligen gjorda uttalande å regeringschefernas vägnar .
stöder kommissionen rådet ?
( en ) fru talman ! när kommissionen i går morse sade att den konstaterar att de åsikter som framförts vara ett gemensamt uttalande av fjorton medlemsstater och att den delar den oro som låg till grund för den åsikten , anser jag att det kan förutsättas att den sedan i går morse och så snart som kommissionen kunde diskutera frågan den haft samma åsikt som de fjorton medlemsstaterna .
tack , kommissionär kinnock .
jag tror att vi upplevt en stor politisk debatt , i nivå med situationen och vad man kunde vänta sig .
tack , kära kolleger .
jag förklarar den aktuella och brådskande debatten avslutad .
tillämpning av försiktighetsprincipen
nästa punkt på föredragningslistan är meddelande från kommissionen om tillämpning av försiktighetsprincipen .
. ( en ) jag vill börja med att säga att jag är glad att få lägga fram detta meddelande om tillämpning av försiktighetsprincipen , och det har författats tillsammans med david byrne och erkki liikanen .
försiktighetsprincipen är inte ett nytt koncept .
den har tillämpats av gemenskapen ganska länge nu på en rad politikområden som miljö , folkhälsa , djur- och växtskydd och den nämns uttryckligen i miljöbestämmelserna i eg-fördraget efter maastricht .
den återfinns även i en rad internationella texter , till exempel rioförklaringen och allra senast i biosäkerhetsprotokollet .
innebörden i försiktighetsprincipen är uppenbar .
den handlar om att vidta åtgärder på ett bestämt politikområde när den vetenskapliga delen inte är klarlagd , men där det finns skälig grund till oro för att de potentiella riskerna är tillräckligt stora för att kräva åtgärder .
tillämpningen av försiktighetsprincipen har emellertid fått en ökad uppmärksamhet under senare år .
händelser som bse och dioxinkrisen har stimulerat till en växande offentlig debatt om vid vilka omständigheter försiktighetsåtgärder är berättigade och nödvändiga .
med hänsyn till detta ökande intresse ansåg därför kommissionen att det skulle vara lämpligt att lägga fram ett meddelande för att fastslå kommissionens ståndpunkt om användningen av försiktighetsprincipen .
det finns två huvudsyften med meddelandet .
dels att förklara på ett tydligt och konsekvent sätt hur kommissionen tillämpar och avser att tillämpa försiktighetsprincipen i sin riskbedömning , dels att fastställa riktlinjer för dess tillämpning baserade på motiverade och konsekventa principer .
vi hoppas också att meddelandet skall bidra till att skapa en bättre allmän förståelse för hur risker skall hanteras och att skingra farhågor om att försiktighetsprincipen skulle kunna användas på ett godtyckligt sätt eller som en förvrängd form för skyddstullar .
kommissionens utgångspunkt för att tillämpa försiktighetsprincipen är behovet att garantera en hög skyddsnivå på områdena , miljö , folkhälsa , djur- och växtskydd .
naturligtvis kan denna målsättning inte användas för att rättfärdiga irrationella eller godtyckliga åtgärder , men det innebär att åtgärder fortfarande kan vidtas även i situationer där vetenskapen är oklar .
medan försiktighetsprincipen inte innebär att man gör politik av vetenskap , vilket några har velat göra gällande , för den oss fram till vägskälet mellan vetenskap och politik .
det inledande beslutet att tillämpa försiktighetsprincipen beror till stor del på den skyddsnivå som eftersträvas och den risknivå som beslutsfattare är beredda att godta för samhället .
den är därför politisk till sin natur .
de åtgärder som senare kan vidtas måste självklart följa de allmänna principer som tillämpas för hantering av risker och riktlinjerna för att tillämpa försiktighetsprincipen är därför den viktigaste delen i dokumentet .
de åtgärder som vidtas skall stå i proportion till den valda skyddsnivån - det vill säga , vi använder inte en hammare för att knäcka en nöt .
de måste vara icke-diskriminerande i sin tillämpning , det vill säga , åtgärder bör inte skilja sig på grundval av geografiskt ursprung .
och de måste överensstämma med redan vidtagna åtgärder .
exempelvis om en produkt har blivit godkänd , bör likartade produkter också godkännas .
åtgärder baseras på en granskning av eventuella fördelar och kostnader för åtgärder eller brist på åtgärd ; det vill säga åtgärderna skall vara kostnadseffektiva och kunna utvärderas mot bakgrund av ny vetenskaplig information och klart fastslå vem som är ansvarig för att lägga fram de vetenskapliga bevis som krävs för en mer djupgående riskbedömning , det är bevisbördan .
alla dessa element skall tillämpas kumulativt .
det är också viktigt att komma ihåg att det finns ett brett urval av åtgärder som kan vidtas vid tillämpning av försiktighetsprincipen .
till exempel ett forskningsprogram , allmänna informationskampanjer , rekommendationer och så vidare .
att tillämpa försiktighetsprincipen medför därför inte automatiskt ett förbud .
det första meddelandet är inte avsett att bli det slutgiltiga ordet i denna fråga . men det är första gången som kommissionen har lagt fram ett strukturerat dokument om principen och dess tillämpning .
genom att fastlägga någorlunda detaljerat hur kommissionen tillämpar och avser att tillämpa försiktighetsprincipen hoppas vi kunna klargöra situationen på gemenskapsnivå och att medverka i den pågående debatten på europeisk och internationell nivå .
herr talman , fru kommissionär ! tack så mycket för förklaringen .
jag har tre mycket korta frågor .
den första frågan : vi har fått vänta mycket länge på ett enhälligt yttrande från kommissionen om försiktighetsprincipen , och tidigare har det över huvud taget inte stått klart om kommissionen talar med en röst .
är det som ni i dag här har lagt fram också den åsikt som era kolleger med ansvar för industri , utrikeshandel , konkurrens och den inre marknaden har ?
ni kommer säkert att säga ja , men jag vill få veta följande av er : känner dessa herrar till vilka konsekvenser det får ?
nästa fråga , fru wallström : när kommer ni att börja att tillämpa detta i lagstiftningen , när det gäller exempelvis kemikalier eller lagstiftning på andra områden ?
den sista frågan : kommer vi att kunna urskilja var detta tillämpats i lagstiftningen ?
det betyder : kommer det att finnas en extra sida i varje förslag som talar om att försiktighetsprincipen har tillämpats och att man kommit fram till detta resultat ?
( en ) tack så mycket , dagmar roth-behrendt , för dessa frågor .
naturligtvis delas detta av hela kommissionen .
detta är ett allmänt meddelande som skrevs av oss tre , david byrne , erkki liikanen och jag själv , men det har godkänts enhälligt i kommissionen i dag .
det fick starkt stöd från övriga kommissionärer och samråd om det har hållits i hela kommissionen .
så vi har verkligen genomarbetat detta dokument och jag är säker på att de alla kan beskriva de riktlinjer och principer som fastslås i detta dokument .
ja , jag kan säga att vi redan använder detta sätt att arbeta med olika , svåra frågor som en ny kemisk strategi till exempel .
jag är också säker på att vi uttryckligen kommer att nämna den när vi arbetar med denna princip .
vi har nyligen haft ett fall där vi använde försiktighetsprincipen när vi måste förbjuda phtalater i mjuka pvc-leksaker och naturligtvis använder vi den på flera olika miljöområden .
den har framför allt använts på miljöområdet , men naturligtvis också när det gäller folkhälsan .
så vi skall försöka vara mycket tydliga om hur och när den skall användas .
herr talman , fru kommissionär ! när det gäller förhållandet mellan vetenskapen å den ena sidan och försiktighetsprincipen å den andra sägs det i meddelandet att det alltid krävs ett politiskt beslut för att använda försiktighetsprincipen när de vetenskapliga bevisen är bristfälliga .
på det sättet lägger man naturligtvis över en hel del makt i händerna på vetenskapen .
man kan undra vilken sorts vetenskapsmän som kommer att lämna den dokumentationen och vad står de för ?
i meddelandet står också att om det finns en tillräckligt stor erkänd minoritet av vetenskapsmän så räcker det för att kunna hänvisa till försiktighetsprincipen .
jag skulle vilja fråga , vad är då definitionen för en erkänd minoritet ?
hur beskriver ni en sådan ?
hur kommer ni fram till en erkänd minoritet ?
när det gäller det politiska beslutet så skulle jag också vilja fråga : vem fattar det politiska beslutet ?
är det rådet ?
i vilken utsträckning kommer parlamentet att kunna delta i det beslutsfattandet ?
vilken funktion har den vetenskapliga kommittén ?
vilken roll kommer inom kort den myndighet för livsmedel som ni skall inrätta att spela ?
avslutningsvis , kommer hela beslutsfattandet att ske på ett öppet och genomblickbart sätt ?
det är mina tre frågor .
( en ) ja , herr talman , det är sant .
det fanns många och svåra frågor och inte alltid kristallklara men jag skall försöka besvara några frågor .
vem vill fatta beslutet , vilka är beslutsfattarna ?
jo , det beror på vilka lagstiftarna är .
detta är en del av riskhantering .
de måste granska exempelvis omsorg om människor i förhållande till en särskild fråga och de måste göra en bedömning mot bakgrund av vad som är känt om vetenskapliga bevis i ett bestämt fall .
men det är sant att det krävs inte uppbackning av en stor majoritet av det vetenskapliga samfundet för att kunna använda försiktighetsprincipen .
den kan tillämpas på basis av bevis från en minoritet eller när vetenskapliga bevis är ofullständiga .
det är naturligtvis där som ni gör en avvägning mellan denna princip som ett politiskt verktyg och vetenskap .
det är inte alltid lätt att beskriva exakt hur denna process fungerar , men det är inte tal om att förändra den vetenskapliga grunden .
vi använder experterna för att få så mycket vetenskaplig information och fakta som möjligt innan vi fattar ett beslut - och det bör också ske i framtiden .
ni måste betrakta denna princip som ett verktyg för riskhantering .
ni måste besluta om ni vill utsätta människor för fara till exempel , eller om ni vill skydda miljön , och ni måste utvärdera de vetenskapliga bevis som finns tillgängliga .
ni måste bedöma allt detta och utvärdera vad vetenskapen visar .
därefter beslutar ni om att vidta en åtgärd eller inte , att göra något eller inte .
således finns det inga svar på alla era frågor , men det förändrar inte det system med forskare som vi använder i dag , eller det system med experter som vi använder i dag .
herr talman ! jag har en fråga som gäller ett konkret och aktuellt fall , i vilket försiktighetsprincipen skulle kunna tillämpas .
det gäller bromerade flamskyddsmedel .
det är så att dessa ämnen nu upptäcks ; det finns ökade koncentrationer av dem i både människor och miljö .
det finns många som hävdar att de medför stora risker , medan andra ifrågasätter hur stora riskerna är med dessa ämnen .
nyligen uppmanade både sverige och danmark i ministerrådet kommissionen att ta ett initiativ för ett förbud mot bromerade flamskyddsmedel .
jag undrar då om ni förbereder ett sådant förbud och om det inte skulle passa väldigt väl in i er syn på själva försiktighetsprincipen att komma med ett sådant initiativ .
herr talman ! tack så mycket , jonas sjöstedt , för denna fråga .
frågan om bromerade flamskyddsmedel är viktig .
den väcktes alldeles nyligen i miljörådet av ett antal ministrar som vill att kommissionen skall titta på vad det finns för underlag och vad som kan behöva göras .
vi är i färd med att se på denna fråga och bedöma vilka kunskaper vi har i dag och vad som är möjligt att göra .
låt mig dock få påminna om att användning av försiktighetsprincipen inte behöver vara samstämmigt med att det skall bli ett förbud , ett totalförbud .
det kan finnas en rad olika åtgärder som kan vidtas .
därför skall det inte omedelbart tolkas som ett förbud .
vad gäller de bromerade flamskyddsmedlen kan det så småningom ändå bli det , men det är viktigt att säga att försiktighetsprincipen tillåter att man använder hela spektrumet av politiska insatser och åtgärder .
denna fråga är aktuell i allra högsta grad .
kommissionen skall göra sitt jobb och titta ordentligt på den innan vi återkommer med en bedömning av vad som behöver göras .
ni framförde att försiktighetsprincipen inte bör användas som ett förtäckt handelshinder .
är denna uppfattning överensstämmande på båda sidor om atlanten ?
jag tror att vi kommer att få problem med i synnerhet hormonbehandlat kött och genetiskt modifierade grödor .
kommer amerikanerna att ha samma uppfattning i denna fråga som vi ?
herr talman ! jag är glad att kunna meddela att vi i montreal precis har skrivit under ett protokoll om biosäkerhet .
där lyckades vi enas i ett internationellt forum om definitionen av försiktighetsprincipen .
jag anser att det är ett genombrott , att vi lyckades avsluta detta protokoll .
jag tror att det kommer att bilda skola för framtida diskussioner om försiktighetsprincipen .
vi kommer att kunna använda detta som ett exempel på hur man skall tolka försiktighetsprincipen .
den är dessutom även accepterad som ett viktigt och verkningsfullt instrument .
jag har två frågor ; jag skall försöka fatta mig väldigt kort .
den första frågan gäller genomförandet av försiktighetsprincipen .
som jag har förstått det , har det varit vissa oklarheter om hur man skall uppfatta detta .
är det så att man först skall göra en riskbedömning där man inkluderar en kostnads- och nyttoanalys , alltså en cost-benefit-analys ?
i så fall blir jag ganska orolig , eftersom det väl var meningen att man inte skall använda en cost-benefit-analys som ett redskap för att avgöra om man skall introducera försiktighetsprincipen , utan försiktighetsprincipen skall komma först .
min andra fråga gäller bevisbördan .
jag minns när margot wallström introducerades som kommissionär i utskottet .
då var hon inne på att man skulle vilja ha en omvänd bevisbörda .
det vill säga att tillverkaren av en produkt skall visa om den är farlig eller inte .
jag vill veta om detta också gäller i det dokument som kommissionen har presenterat nu .
tack så mycket , inger schörling .
detta är två viktiga frågor .
det är bra att jag får tillfälle att klargöra dem .
nej , man måste inte börja med att göra en cost-benefit-analys , utan detta skall baseras på en bedömning av vad vi vet , vad vetenskapen kan berätta för oss och hur vi skall se på det jämfört med de risker som vi bedömer finns för miljön eller för hälsan hos människor och djur .
däremot när man har bestämt sig för att vidta en viss åtgärd , då bör man välja en kostnadseffektiv åtgärd , så att man faktiskt inte tar till åtgärder som är helt orimliga när det gäller effektivitet .
det är alltså inte så att man måste börja med en cost-benefit-analys .
den andra frågan rör den omvända bevisbördan .
det är alldeles riktigt att vi behöver tillämpa det i vissa fall .
jag har använt exemplet kemikaliestrategin som ett bra exempel på ett område där vi behöver göra detta .
då handlar det emellertid om det sakområdet , medan man kan säga att detta meddelande om försiktighetsprincipen är horisontellt ; det gäller alla olika specifika politiska sakområden .
därför diskuteras inte speciellt i detta sammanhang en omvänd bevisbörda eller hur bevisbördan skall se ut , utan det handlar i stället om det politiska beslutsfattandet och grunderna för detta .
det är dock alldeles riktigt att vi t.ex. när det gäller kemikalier måste se till att vi får en omvänd bevisbörda .
herr talman ! jag anser att försiktighetsprincipen för att fungera måste tillämpas ganska radikalt , för annars förlorar vi oss i tolkningarnas irrgångar .
låt mig ge ett exempel : det visar sig att en antikryptogam gör så att det föds blinda barn , medlet är med andra ord teratogent .
ok , detta är en antikryptogam , ett antimögelmedel .
den teratogena effekten har påvisats av ett enda engelskt laboratorium , kanske det enda laboratorium som har gjort några undersökningar .
jag anser då att försiktighetsprincipen , med tanke på att det rör sig om ett så allvarligt hot mot hälsan , kräver att produkten omedelbart skall förbjudas , så som till exempel nya zeeland har gjort .
låt mig alltså ställa den här frågan : när människors hälsa står på spel , eller man riskerar allvarliga hälsoeffekter , skall man då kanske göra en kostnads / intäktsanalys ?
den kostnad som ett blint barn innebär är enligt mitt förmenande alltför hög , det finns inga vinster som kan uppväga den .
jag vill därför veta om försiktighetsprincipen i det här fallet , så som ni tolkar den , fru kommissionär , förutsätter att produkten under alla omständigheter skall tas ur marknaden till dess att bevis om motsatsen har framlagts av andra laboratorier .
herr talman ! jag är den första att önska att vi kan tillämpa försiktighetsprincipen på ett sådant sätt att det upplevs som radikalt till skydd för människors hälsa och för miljön .
det är klart att jag inte kan ta ställning till det speciella fall och den speciella produkt som nämns här , men jag skall direkt gå tillbaka och se vilken information jag kan få fram om just detta fall .
sanningen är ju att väldigt många medlemsstater , förvisso också andra nationer , har vidtagit åtgärder för att skydda sin befolknings hälsa på ett sådant sätt att man har använt försiktighetsprincipen , även om man inte alltid har kallat det så .
det är naturligtvis så att det inte i första hand är frågan om en kostnad ; det kan nämligen bli en enorm kostnad för samhället om man undviker att vidta en viss åtgärd .
det får inte heller vara så att man sitter och räknar vad ett människoliv kostar gentemot att vidta en åtgärd .
jag tycker dock att det är alldeles självklart att när det så småningom är dags att besluta sig för en åtgärd , är det ofta så att man har många olika handlingsalternativ .
då skall man titta på vad som ger bäst resultat .
jag kan inte låta bli att berätta om ett tillfälle när detta uttryck användes av personer som man kanske inte alls skulle kunna tänka sig använda ordet kostnadseffektiv , nämligen vid ett besök i afrika .
på ett hospice för aidspatienter träffade jag två irländska , katolska nunnor som skötte om döende aidspatienter .
de var de första att säga att vi måste varje dag tänka på att göra det som är mest kostnadseffektivt , därför att det måste räcka till våra stackars patienter här ; vi måste vara mycket noga med hur vi använder resurserna .
jag menar att vi kan lära oss något av detta .
vi måste ju alltid se till att vi använder våra resurser på effektivaste sätt och så att de kommer till hjälp på bredast möjliga sätt .
det är alltså inte korrekt att man först måste börja med någon sorts cost-benefit-analys , vilket också förklaras i detta meddelande .
man skall titta på vad vetenskapen erbjuder för kunskaper , och man skall använda detta som ett viktigt politiskt instrument för att skydda miljön och människors hälsa .
herr talman ! det är en sällsynt nåd att få en andra möjlighet att ställa en fråga !
fru kommissionär , jag vill än en gång komma tillbaka till min första fråga , som kanske lät skämtsam , när jag frågade efter de andra kommissionärerna .
ni besvarade den också så som jag visste att ni skulle göra .
jag skulle vilja knyta samman den med något som goodwill frågade , nämligen med vårt förhållande mellan försiktighetsprincipen och världen utanför europeiska unionen .
jag frågar ju inte detta utan orsak .
ni har med all rätt sagt att försiktighetsprincipen är nödvändig just när vetenskapen ännu inte har några bevis .
hur skall vi se till att vi inte alltid blir möjliga att angripa , t.ex. av våra partner i usa - och då räcker inte bio safety-protokollet till ?
hur skall vi se till att inte industripolitikerna och utrikeshandelspolitikerna sparkar undan benen för er på samma sätt som de tidigare alltid gjorde med era företrädare ?
det är just det som det handlar om , annars behöver vi här inte tala om försiktighetsprincipen , fru kommissionär !
herr talman ! jag tycker att det är väldigt viktigt att visa på de riktlinjer som finns för användande av försiktighetsprincipen i detta meddelande som ett sätt att tillbakavisa påståendena om att vi alltid vill använda detta av protektionistiska anledningar .
jag är säker på att vi kommer att få fler konflikter med t.ex. usa .
vi skall inte vara naiva och tro något annat .
ända sedan vi skrev under detta protokoll i montreal , har vi emellertid ett internationellt erkännande och en gemensam definition inskriven i ett protokoll som handlar om miljö , hälsa och handel .
det utgör därför ett gott exempel .
vi skall inte tro något annat än att det kan dyka upp konflikter även i fortsättningen , men nu kan vi visa att vi inte använder försiktighetsprincipen godtyckligt .
vi har nu ett antal riktlinjer för detta , och vi har ett starkt stöd hos våra respektive befolkningar för att använda försiktighetsprincipen , vilket tydligt fastläggs i detta meddelande .
den uppmärksamhet som ägnats åt den politiska försiktighetsprinipen har lett till att vi har diskuterat frågan i ungefär två timmar och nu anses den frågan så att säga ligga utanför den normala rutinen , även om , som vi har kunnat konstatera av de inlägg vi har hört i dag , från frågorna och svaren , det är en fråga som man fäster stor vikt vid .
nästa punkt på föredragningslistan är betänkande ( a5-0018 / 2000 ) av dimitrakopoulos och leinen för utskottet för konstitutionella frågor om sammankallandet av regeringskonferensen ( 14094 / 1999 - c5-0341 / 1999 - 1999 / 0825 ( cns ) ) .
( el ) herr talman ! jag skall till att börja med tacka det portugisiska ordförandeskapet och kommissionen för alla de mycket nyttiga kontakter som vi har haft under denna tid .
tillåt mig även att än en gång tacka min medföredragande , leinen , för allt vårt samarbete .
herr talman , kära kolleger ! den regeringskonferens som skall starta är viktig , både rent allmänt , men särskilt med tanke på den förestående utvidgningen .
vid denna skall den struktur och den metod som skall ligga till grund för europas funktion i det 21 : a århundradet utarbetas .
för att europeiska unionen i framtiden skall kunna fungera effektivare , mer demokratiskt och med full öppenhet , är det uppenbart att det krävs en omfattande och grundlig reform av europeiska unionens institutioner liksom av deras arbetsmetoder .
av avgörande betydelse för att denna reform skall lyckas är den dagordning som skall ligga till grund för arbetet på regeringskonferensen .
av besluten från toppmötet i helsingfors framgår att den dagordning som man där kom överens om inte är tillfredsställande , och att den inte garanterar de nödvändiga och påtagliga förändringar som är ett måste för att skapa ett europa som fungerar bättre , är effektivare , mer demokratiskt och mer öppet .
och detta på grund av att den är begränsad till endast de tre frågor som på ett lösryckt sätt berör strukturen och funktionen hos endast två av europeiska unionens institutioner .
jag skall inte upprepa det , för ni känner väl till det allihop .
detta mitt konstaterande berättigas dels av det ständiga kravet från de europeiska medborgarna , som till och från är mycket kraftigt , dels av de enorma dimensionerna på det projekt som europeiska unionen redan har gett sig in i , utvidgningen .
mot denna bakgrund är det inte möjligt att man i dagordningen för den nya regeringskonferensen inte inbegriper frågor som , om de får en lösning , skulle säkerställa en smidig funktion för alla - inte bara vissa - av europeiska unionens institutioner .
liksom det inte heller är möjligt att man i dagordningen inte inbegriper frågor som dagligen berör och som därför är mycket påtagliga för den europeiska medborgaren .
herr talman , kära kolleger ! europaparlamentet har under sina många diskussioner och i de betänkanden som har lagts fram till dags dato öppet varit för att sammankalla en regeringskonferens .
jag begär emellertid att man på denna parallellt skall ta upp både frågor som förbättrar och fullbordar reformen av - och jag upprepar det - alla institutioner och frågor som direkt berör och intresserar de europeiska medborgarna . som till exempel hälsa , energi , kultur , transport och till och med turism .
vad gäller frågan om dagordningen till slut kommer att utvidgas eller inte , är den å ena sidan fortfarande under diskussion . och här vill jag verkligen prisa det sätt på vilket det portugisiska ordförandeskapet , som vid upprepade tillfällen inför europaparlamentet har förbundit sig att arbeta i den riktningen , har uppträtt politiskt .
å andra sidan får en ökning eller ett bevarande av antalet frågor inte under några omständigheter leda till att den betydelse som varje medlemsland tillskriver regeringskonferensen minskar .
och detta av den anledningen att den institutionella ram som skall ligga till grund för europa i framtiden är en grundläggande princip för den europeiska integreringen och följaktligen en fråga av högsta nationella betydelse för varje land som är medlem i unionen .
herr talman , kära kolleger ! med detta som bakgrund uppmanar jag kammaren att godkänna det yttrande som jag och leinen har lagt fram , så att regeringskonferensens arbete kan komma igång den 14 februari och så att våra två företrädare på denna , brok och tsatsos , kan gå framåt med europaparlamentets samtycke i det svåra arbete som de har framför sig .
samma sak gäller även för europeiska kommissionen , och jag vill , återigen , tacka kommissionär barnier för hans kontakter med europaparlamentet och för de mycket konstruktiva förslag som han har lagt fram för oss .
herr talman ! europeiska folkpartiets grupp ( kristdemokrater ) och europademokrater var inte nöjda med resultatet från europeiska rådets möte i helsingfors .
vi ansåg att dagordningen var för begränsad , för vår grupp utgick från fördragets logik , närmare bestämt från protokollet om unionens institutioner .
i helsingfors kom regeringarna överens om att en minimireform är tillräcklig , så länge europeiska unionen består av mindre än 21 stater ; dessutom krävs det en djupgående reform .
samtidigt godkände europeiska rådet i helsingfors en utvidgning med 13 nya medlemsstater .
det finns således en motsägelse i att påbörja anslutningsförhandlingarna med 13 samtidigt som man vill ha en minimireform .
vi tillämpar fördragets logik och vill att dagordningen för nästa regeringskonferens skall rymma en mer djupgående reform av unionen .
det är anledningen , herr talman , till att vi håller denna debatt i parlamentet i dag , eftersom vi inte vill skjuta upp inledandet av konferensen .
rent teoretiskt hade vi kunnat göra det .
vi hade kunnat rösta den sjuttonde den här månaden , och då hade inte konferensen kunnat börja den fjortonde .
men det ville vi inte göra , för vi vill ge regeringarna och kandidatländerna en tydlig politisk signal om att vi önskar genomdriva denna reform just för att underlätta en utvidgning .
herr talman , jag är glad över att kunna framföra detta till det portugisiska ordförandeskapet , för de har vunnit ett gott anseende här i parlamentet .
det portugisiska ordförandeskapet delar många av parlamentets ambitioner , och man har lovat att göra vad man kan för att regeringskonferensens dagordning skall fyllas på med andra frågor som är av största vikt .
och jag vill dessutom påpeka , herr talman , att europaparlamentets ambitioner inte är ambitioner för parlamentets egen räkning .
europaparlamentet kommer hur som helst att stärkas politiskt av det fördrag som regeringskonferensen resulterar i .
anledningen till detta är mycket enkel : under regeringskonferensen kommer man , i enlighet med överenskommelsen i helsingfors , att ta ställning till vilka av de frågor som hittills har avgjorts med enhällighet som skall avgöras med kvalificerad majoritet .
det innebär att antalet frågor som avgörs med kvalificerad majoritet kommer att öka .
och det framgår redan av gemenskapens regelverk att de lagstiftningsfrågor som avgörs med kvalificerad majoritet även skall vara föremål för parlamentets medbeslutande .
därför innebär en ökning av den kvalificerade majoriteten en ökning av parlamentets medbeslutande .
däremot skulle parlamentet inte uppfylla sin roll som en supranationell europeisk institution om det inte tänkte på unionens politiska utformning .
det är det vi ägnar oss åt nu .
vi anser att unionens politiska utformning förutsätter att även andra frågor behandlas .
bland annat sådana som handlar om införandet i fördraget av säkerhets- och försvarsfrågor , frågor vars betydelse har ökat markant den senaste tiden och därför bör införlivas i fördraget .
förvisso även stadgan om de grundläggande rättigheterna i europeiska unionen , vars utformning påbörjades i går , och jag tror att man gripit sig an den uppgiften på ett mycket positivt sätt .
vi kommer i stor utsträckning att verka för att européerna skall bli medvetna om fördelarna med att vara europé och att en europeisk medborgare har vissa grundläggande rättigheter som är knutna till unionens institutioner .
de förslag , herr talman , som vi konkretiserar i ett annat betänkande , utgör tillsammans med kommissionens förslag ett utmärkt dokument som - vilket jag nu har nöjet att få säga till herr barnier - således kommer att vara ett underlag till regeringskonferensen .
det får vi tala mer om en annan dag .
i dag måste vi ge klartecken till sammankallandet av denna konferens , och europeiska folkpartiets grupp , herr talman , är beredd att ge klartecken .
herr talman ! å socialistgruppens vägnar kan jag framföra att vi kommer att stödja det förslag till yttrande som lagts fram av föredragandena för utskottet för konstitutionella frågor .
vi avger ett positivt yttrande om att sammankalla regeringskonferensen helt enkelt därför att vi är mycket imponerade av det portugisiska ordförandeskapet som har gått med på vår begäran om att dagordningen för regeringskonferensen utvidgas .
resterna från amsterdam är inte ett bra uttryck eftersom de är mycket viktiga frågor i sig själva .
låt oss kalla dem de tre första punkterna för regeringskonferensen .
dessa tre första punkter är mycket viktiga , men detta är frågor som diskuterades noga av våra medlemsstater under den senaste regeringskonferensen .
de kom inte helt fram till en slutsats om dem men det krävs verkligen inte nio månader av ytterligare granskning av dem .
de kräver en politisk överenskommelse .
det är mer en fråga om nio minuter , kanske nio timmar om det är svårlöst , inlåsta tillsammans i ett rum för att nå en lösning om dessa frågor , inte nio månader .
under dessa omständigheter skulle det vara dumt att inte utvidga dagordningen .
det finns andra frågor som borde vara givande att granska framför allt före en så stor utvidgning av unionen med så många nya länder .
ingen begär att det ska vara julklappsstämning .
ingen begär en regeringskonferens i stil med maastricht med hundra eller fler punkter att diskutera .
men det finns sex , sju , åtta , kanske nio punkter som det skulle vara mycket lämpligt och nyttigt att få en lösning på .
det finns tid .
kom ihåg regeringskonferensen som ledde fram till europeiska enhetsakten .
den pågick bara fem månader .
den regeringskonferens som ledde fram till det enorma maastrichtfördraget pågick ett år .
enbart konferensen om amsterdamfördraget pågick i ett och ett halvt år och det berodde på att alla visste att man måste vänta på resultaten av det brittiska valet om man skulle få något resultat från den regeringskonferensen , så det var av en annan orsak .
ett år är tillräcklig tid för att lösa en stort antal frågor , och det borde utan tvivel vara tillräcklig tid för att lösa de få avgörande frågor som vi önskar lägga till på dagordningen .
jag är glad att kommissionen delar vår åsikt .
kommissionen har just offentliggjort sitt yttrande och den har gjort exakt det som parlamentet begärde av den - att lägga fram ett fullständigt och samlat förslag med verkliga förslag till fördragsartiklar .
jag tackar kommissionen för detta även om jag naturligtvis inte är överens med allt det som kommissionen framförde .
jag anser att det finns några brister i det som den presenterade .
hur som helst har kommissionen tillhandahållit en tjänst och jag uppskattar att kommissionär barnier som finns här bland oss i dag för att han gjorde detta .
den har för allmänheten presenterat några av de avgörande frågor som vi måste lösa under denna regeringskonferens .
det är alltsammans bara bra .
parlamentet , rådets ordförandeskap och kommissionen drar åt samma håll för att få en bredare dagordning .
jag önskar er all framgång , rådets ordförande , för att se till att europeiska rådet godkänner denna dagordning och att på alla hjärtans dag när ni inleder regeringskonferensen det kommer att ske under gynnsamma omständigheter och att ni kommer att kunna slutföra den på ett bra sätt , även när det franska ordförandeskapet tar över i slutet av detta år .
vi skall inte längre oroa oss över att dagordningen för regeringskonferensen skall bli begränsad .
det är en av de politiska slutsatserna som vi måste dra från det allvarliga beslutet av 14 medlemsstater i går att i verkligheten frysa våra förbindelser med en partner .
det gör det omöjligt för dessa samma medlemsstater att vid regeringskonferensen misslyckas med att ge en effektiv mening vad gäller skydd och främjande av grundläggande fri- och rättigheter .
det är redan konstigt att inom det konvent som tar fram förslag till stadgan se företrädare från några medlemsstater , särskilt storbritannien och frankrike , försöka argumentera att en obligatorisk stadga på något sätt skulle vara en kränkning av nationellt självbestämmande .
det är viktigt att regeringskonferensen förbereder hur införandet av en ordning för grundläggande fri- och rättigheter inom fördraget godkänns .
en del av detta är att förbättra medborgarnas möjlighet att väcka talan vid domstol .
ett annat sätt är att själva unionen undertecknar europakonventionen .
ett annat sätt är utan tvivel att nationella parlament och nationella politiska partier finna en kraftfullare roll som de kan spela inom europeiska unionens verksamhet och att dela ansvaret för att skapa europeisk parlamentarisk demokrati .
min grupp välkomnar absolut regeringskonferensen och kommer att medverka i denna fördragsreform i största möjliga grad .
herr talman ! gruppen de gröna / europeiska fria alliansen anser att europaparlamentets beslut att skyndsamt yttra sig om regeringskonferensen neutraliserar den politiska betydelsen av uppmaningen till rådet och gör den , i slutändan , ganska ointressant .
vi hade hellre velat få en tydligare uppfattning om dagordningen , något större säkerhet vad gäller metoden , innan vi avger vårt yttrande , och vi uppskattar inte den bristande respekt som det portugisiska ordförandeskapet visade europaparlamentet genom att bestämma att regeringskonferensen skulle börja på alla hjärtans dag , den första dagen under sammanträdesperioden i strasbourg .
jag tror dessutom att eftersom detta är ett ganska viktigt yttrande , så kan vi också rösta för det och jag tror att majoriteten i vår grupp kommer att rösta för det .
man jag vill ändå understryka att det är ganska grymt att se hur litet intresse denna reform väcker .
händelserna i österrike visar på ett mycket tydligt sätt behovet av en reform , en struktur för den europeiska demokratin , för att bestämma de principer som samtliga medlemsstater skall ansluta sig till .
det smärtar också att tänka sig att initiativet gentemot österrike i verkligheten är frukten av en överenskommelse mellan regeringar och att europeiska unionen och dess institutioner inte hade möjligheter eller den gemensamma kraften att agera för att förhindra utvecklingen och leda in den på andra banor .
jag tror att detta är något som vi måste reagera mot , detta måste vi göra under regeringskonferensen och jag hoppas verkligen att europaparlamentet inte med det här yttrandet , som avgivits med sådan ovilja , helt har uttömt sin förmåga att utöva påtryckningar på rådet och medlemsstaterna för att denna regeringskonferens inte bara skall bli en rent teknisk övning utan väcker den entusiasm som vi fick se spår av i detta parlament för några timmar sedan .
herr talman , herr rådsordförande , herr kommissionär , ärade kolleger ! jag anser att man inte tillräckligt ofta och ljudligt kan säga att den föredragningslista som rådet har fastställt för regeringskonferensen är politiskt fullständigt oacceptabel , och jag vill tillfoga att jag anser att den rent av är skamlig .
vi befinner oss nämligen i en historisk situation , där man förhandlar respektive kommer att ta upp förhandlingar med 12 stater , och nu befinner vi oss gemensamt i en situation där det inom överskådlig tid kan bli verklighet att europa växer samman .
men hur skall då unionen kunna utvidgas , om man inte nu - alltså före utvidgningen - ser till att man har effektiva verktyg ?
därför är vi som grupp positiva till regeringskonferensen .
vi anser att den är absolut nödvändig och brådskande och vi hoppas att den i själva verket skall åstadkomma resultat som möjliggör en snar utvidgning av europeiska unionen .
min grupp , herr rådsordförande , har med tillfredsställelse noterat att rådets ordförandeskap inte är tillfreds med den nuvarande situationen .
därför kan ni vara säkra på att även gruppen europeiska enade vänstern / nordisk grön vänster kommer att arbeta för att unionen äntligen skall göra sina hemläxor .
det handlar om varken mer eller mindre än europas framtid , och det handlar framför allt om ett europa som medborgarna faktiskt uppfattar som sitt eget , eftersom de kan vara med och utforma det , och eftersom de bekymmer och trångmål , problem och frågor som de dagligen möter också tas på allvar i politiken .
de slutna dörrarnas politik , samråden i den stilla kammaren , allt detta måste en gång för alla förpassas till det förflutna .
därför krävs det öppenhet .
jag anser att ni som ordförandeskap bör se till att tåget inte fortsätter att gå som hittills , och att människorna inte blir stående kvar på perrongen som fördragsanalfabeter .
vi anser att det är absolut nödvändigt att man inte bara gör allt för att ge medborgarna omfattande information om vad som sker vid regeringskonferensen och resultaten av den , utan de måste snarare integreras direkt i hela reformprocessen .
vi anser också att de politiska beslutsfattarna äntligen måste hoppa över sin skugga och efter regeringskonferensen fråga medborgarna i folkomröstningar om de är införstådda med hur deras europa kommer att utvecklas i framtiden .
på så vis skulle vi faktiskt få ett medborgarnas europa , och vi skulle faktiskt få en helt ny kvalitet med demokratisk legitimitet för unionen .
jag vill klart och tydligt ta upp en annan central demokratifråga .
som ledamot av den församling , som nu har påbörjat sitt arbete på stadgan för de grundläggande rättigheterna , vill jag klart säga : för mig och min grupp räcker det inte med att högtidligt förkunna stadgan .
vad kommer väl medborgarna att säga när man högtidligt förkunnar rättigheter för dem , medan de inte som individer kan överklaga något ?
nej , jag tror att det bara skulle fördjupa unionens trovärdighetskris ännu mer .
det dåliga valdeltagandet vid europavalen bör verkligen vara en tillräcklig larmsignal för alla .
det vi behöver är synliga rättigheter för var och en , stadgan om de grundläggande rättigheterna måste blir bindande rätt för alla människor som bor i unionen , för alla dess medborgare .
detta är det mål som vi för medborgarnas skull gemensamt bör arbeta för , och jag förväntar mig av regeringskonferensen att beslutet från köln i denna fråga revideras vid årets slut .
naturligtvis handlar det också om att man har effektiva beslut och fungerande institutioner i en union med 27 och fler medlemsstater .
med enbart en liten minireform , som rådet har bestämt sig för , kommer det inte att lyckas , och därför bör alla institutioner prövas .
vi behöver modiga förändringar , och därvid måste vi samtidigt se till att man ägnar största uppmärksamhet åt jämställdheten mellan de stora och de små staterna .
detta vill jag särskilt betona som ledamot från ett stort medlemsland .
jag tackar kommissionen för de förslag den har lagt fram , och jag är säker på att vi här kommer att få omfattande diskussioner med medborgarna även i europaparlamentet om alla de frågor som de har framkastat .
jag vill också ta upp en sista fråga .
i parlamentets yttrande krävs det uttryckligen ändringar av fördraget när det gäller den ekonomiska politiken .
i själva verket är det så att globaliseringen av samhällsekonomin , men framför allt införandet av euron och den stabilitetspakt som är förbunden därmed , gör det nödvändigt att inte bara fråga efter bakgrunden till beslutsprocesserna .
det som framför allt krävs är modet att kritiskt granska unionens hittillsvarande politik .
det handlar om ett socialt rättvist europa .
ett socialt rättvist europa är oförändrat högaktuellt , ty det handlar i första hand om att målinriktat ställa kampen mot massarbetslösheten och fattigdomen i centrum för unionens politik .
hit hör därför också , enligt min åsikt , modet att ändra artikel 4 i eg-fördraget , som unionen på klassiskt nyliberalt vis definierar som en öppen marknadsekonomi med fri konkurrens , och dit hör enligt min åsikt även artikel 105 i eg-fördraget , ty europeiska centralbanken måste äntligen få ett i fördraget fastslaget politiskt uppdrag att med sin penningpolitik främja hållbar tillväxt och sysselsättning .
herr talman , kära kolleger ! jag talar som företrädare för de italienska radikala ledamöterna och jag skulle vilja säga till rådets ordförande att han förmodligen har kunnat konstatera vad som är parlamentets uppgift .
det är knappast en slump att det sista inlägget var det enda som han instämde i helhjärtat - jag säger detta utan att på minsta sätt ironisera över den position , som är fullständigt respektabel , som berthu och hans grupp har intagit - men det är ingen slump att europeiska rådets beslut stöds av dem som egentligen befinner sig i detta parlament enbart för att de är motståndare till - något som är fullständigt respektabelt - en ytterligare integration i europa .
detta är det budskap som parlamentet skickar till rådet .
jag hoppas att det portugisiska ordförandeskapet - och som även jag vill gratulera - kan överbringa detta parlaments budskap och blir de som bär fram resultatet av vårt kompromissarbete till st .
valentins altare , men under alla omständigheter kommer vi i morgon att yttra oss negativt om dagordningen för regeringskonferensen .
det här budskapet måste bli mycket tydligt : det är så vi tolkar den röst som vi avger i morgon .
vi avger ett yttrande - som är tekniskt och juridiskt nödvändigt - för att sammankalla regeringskonferensen den 14 februari , men vi yttrar oss negativt om innehållet .
det räcker att betänka de faktiska omständigheterna : vi såg österrike för ett tag sedan , men vi kan också se på aktiebörserna , herr talman : när , på ett år , det stora europrojektet kan förlora 16 procent gentemot dollarn så borde kanske inte en regering , men väl en god familjefader , fråga sig om man kan säga till medborgarna att det enda man kan förhandla om är antalet europeiska kommissionärer eller andra frågor av samma typ .
det är uppenbart att målet måste vara ambitiösare .
vi radikala har lagt fram ändringsförslag som vi kommer att underställa kammaren , för att skärpa texten , för att till exempel begära det som borde vara ett minimum - om man nu skall tala om artikel 6 och 7 - dvs. att den europeiska konstitutionen även skall utformas av europaparlamentet , att man föreslår att ändringarna i fördraget skall godkännas av europaparlamentet .
vi vet att det även finns andra frågor : till exempel har många kolleger , tillsammans med oss , skrivit under frågan om var institutionerna skall vara belägna , en fråga som vi tycker borde utgöra en del av de diskussioner som förs under regeringskonferensen .
låt mig avslutningsvis hoppas att det budskap som vi ger i morgon blir ett kraftfullt budskap , för en gångs skull betydelsefullt , och att man verkligen , även tack vare de ansträngningar som det portugisiska ordförandeskapet gjort , kan revidera denna dagordning , för annars tror jag verkligen att detta är ett tillfälle som går förlorat , inte bara för ögonblicket , utan för många år framåt .
herr talman ! kommissionens ordförande var inte helt ärlig när han i förra veckan uttalade sig om regeringskonferensen .
han sade att det fortfarande skulle finnas enhällighet i sociala frågor , men i kommissionens förslag vill man ju uttryckligen ha majoritetsbeslut i socialförsäkringsfrågor och frågor som rör de skatter som har samband med den inre marknaden , och det betyder att huvuddelen av de sociala systemen i medlemsstaterna skall kunna ändras av en majoritet i bryssel , även om en enhällig fransk nationalförsamling , ett enhälligt brittiskt underhus och en enhällig nederländsk andrakammare är emot det .
man går här in i folkstyrets hjärta rörande fördelningspolitiken och medborgarnas sociala villkor , som är det man vill påverka när man går till val .
detta skall vi inte längre kunna bestämma över som väljare . detta skall vi inte längre kunna ändra på valdagen .
bryssel vet bättre .
prodi bebådade också större öppenhet , men hans förslag till förordning innebär en direkt bakåtsträvande utveckling och det är inte bara min , utan också europeiska ombudsmannens uppfattning .
i dag är kommissionen skyldig att individuellt väga sekretesshänsynen mot medborgarnas krav och förväntningar rörande öppenhet , och om kommissionens förordning antas kommer kommissionen att ha att utestänga en rad dokumentkategorier , utan att genomföra en konkret bedömning .
man vill också skapa rättsliga krav på sekretess och sekretessbelägga dokument som i dag är offentliga i en rad medlemsstater .
under titeln &quot; utveckling för öppenhet &quot; gör man att en rad dokument inte blir tillgängliga för allmänheten .
det är mycket orwellskt .
jag vill be prodi att aldrig mer kommentera ett förslag här i kammaren , som inte samtidigt finns tillgängligt för allmänhetens kritiska kontroll .
prodi talade i positiva ordalag om ett förslag som annars hade fått kritik , då det i det nya förslaget till förordning framställs som ett framsteg att man nu skall skapa insyn i alla dokument som finns hos kommissionen , men efteråt kommer en lång , lång lista över undantag , och det finns rättsliga krav på sekretess rörande dessa undantag .
i den franska texten står det &quot; refuse &quot; , i den engelska &quot; shall &quot; , vilket innebär att kommissionen skall hemlighålla uppgifter som i dag är offentliga i t.ex. mitt hemland .
det finns också en gummiparagraf om förhandlingarnas och institutionernas effektivitet , som kan användas till vad som helst , det är därför ...
( talmannen avbryter talaren . ) .
herr talman , kolleger ! efter det portugisiska ordförandeskapets framställning har jag en känsla av att man tar itu med denna regeringskonferens med väl övervägda tankar och ett stort mått av öppenhet .
som europaparlament kommer vi att utnyttja dessa möjligheter för att där på lämpligt sätt lägga fram våra frågor .
kommissionens hittillsvarande förberedelser går åt rätt håll , även om de också enligt europaparlamentets resolutioner inte går tillräckligt långt .
det kommer ju också att diskuteras senare .
det som är avgörande för denna regeringskonferens är att det uppnås en treklang , nämligen handlingsförmåga , demokratisk legitimitet och öppenhet .
endast om dessa tre saker finns för handen , får vi till slut en acceptans från medborgarna .
handlingskraften skall naturligtvis skapas för att det skall vara möjligt för europeiska unionen att utvidgas .
när vi i denna kammare i dag tidigare förde en annan debatt , så är det ett viktigt tecken för detta .
vi måste också vara handlingskraftiga i en europeisk union , om det någon gång skulle hända att en regering skulle utöva en totalblockad .
det är ett viktigt tecken på att majoritetsbeslutet är en avgörande förutsättning för att europeiska unionen skall kunna arbeta i alla sammanhang .
detta är särskilt viktigt i samband med utvidgningen , när det gäller lagstiftning , och när det gäller fördrag som för med sig ändringar av lagstiftningen .
här vill vi naturligtvis också bygga ut motsvarande rättigheter för europaparlamentet .
därvid kommer vi som europaparlament också att agera när det gäller emu , ty på detta område finns det inte någon tillräcklig kontroll .
finansministrarna uppträder i ekofin-rådet och med de 11 staterna i euro-rådet som om det vore ett evenemang mellan regeringar , vilket inte är acceptabelt .
i motsats till kaufmann är jag inte positiv till att utvidga kontrollen av europeiska centralbanken , eftersom jag är för europeiska centralbankens oberoende .
men politiskt sett måste kontrollen åstadkommas på lämpligt sätt .
det gäller också att återställa trojkan kommissionen , rådet och parlamentet i fråga om utrikes- och säkerhetspolitiken , där hittills allt har skötts alltför mycket av rådet , och särskilt de primitiva krisstyrningsåtgärderna , där ansvaret ligger enbart hos kommissionen .
allt detta har inte tagits med i detta helhetskoncept i tillräcklig omfattning .
vi måste granska om det är nödvändigt med ändringar här inom ramen för regeringskonferensen .
rådets portugisiska ordförandeskap har sagt ja till att arrangera överläggningar om detta , för att möjligen få en utvidgning av mandatet .
jag vill också hänvisa till en annan viktig punkt .
de diskussioner vi i dessa dagar för om exempelvis en regering i ett land i europa , visar ändå att vi måste fastslå europeiska unionens intellektuella , moraliska , rättsstatliga inriktning med en gemenskaps- och allmännyttig orientering , och att rättsligt bindande grundläggande rättigheter även av den anledningen måste införas i fördraget , eftersom detta kommer att vara en avgörande stabiliserande faktor .
jag ber dem som i detta avseende hittills har varit mycket återhållsamma , att överväga om det nu inte är rätt ögonblick att också inse detta sammanhang och kanske ha det mod som krävs , så att vi på lämpligt sätt kan komma vidare med de grundläggande rättigheterna .
europeiska unionen behöver knappast några nya instrument , inga nya befogenheter .
det den behöver är instrument för att kunna utnyttja sina befogenheter .
av den anledningen måste vi se till att instrumenten kan fungera så att vi i medborgarnas namn kan utföra de uppgifter , som vi formellt redan har ålagts i fördraget .
jag tror att denna regeringskonferens särskilt bör koncentrera sina ansträngningar på detta .
om vi lyckas uppnå några framsteg här , då kan vi också se fram emot den historiska uppgiften att utvidga europeiska unionen .
det måste vara den avgörande punkten .
ärade ordförandeskap i rådet , jag är övertygad om att det kommer att utformas på ett positivt sätt under er ledning .
ni har säkert , efter att ha lyssnat på de olika inläggen förstått hur uppfattningen att vi skall visa det portugisiska ordförandeskapet förtroende , att vi inte skall öka dess svårigheter genom att skjuta regeringskonferensen på framtiden , har segrat i utskottet för konstitutionella frågor , och även när det gäller ordförandena för de olika politiska grupperna i parlamentet .
jag kan försäkra er att det inte var lätt att lyckas med detta i förra veckan i det utskott som jag leder , men vi har nu definitivt beslutat att satsa på det portugisiska ordförandeskapet , och det är en satsning som vi verkligen hoppas kommer att gå hem .
ni talade om era resor mellan olika huvudstäder och ni berättade om de svårigheter som vissa regeringar har att skapa enighet i sina länder och därmed också i sina respektive parlament .
låt mig påpeka för er att i går genomförde vi en som jag tycker mycket intressant diskussion och dialog med företrädarna för de 15 olika nationella parlamenten , som var närvarande med kvalificerade och engagerade delegationer .
det handlade inte om att komma fram till några slutsatser - det var inte möjligt att dra några sådana - men diskussionerna var utan tvekan mycket uppmuntrande .
jag anser att vi måste vara försiktiga , och verkligen vara övertygade om att de olika nationella regeringarna faktiskt försöker övertala sina respektive parlament att ratificera lösningar som motsvarar behovet att utöka unionen och att inte ta skydd bakom motståndet från sina respektive parlament för att inte underteckna de slutsatser som krävs vid regeringskonferensen .
vi kommer under alla omständigheter att förstärka vårt samarbete , vår dialog med de nationella parlamenten under hela den tid som regeringskonferensen pågår .
i går diskuterade man även inom kommissionen - här företrädd av kommissionär barnier - som också avgav sitt yttrande .
man uppskattade ansträngningarna även om man , när det gäller förslagen , uttryckte avvikande åsikter , i likhet med vad även ni har gjort , herr rådsordförande , om jag inte misstar mig .
det som måste understrykas är det faktum att även i går var många medvetna om risken att utvidgningen leder till att den ursprungliga idén att bygga upp ett politiskt europa kan komma att ifrågasättas , en risk som för övrigt påpekades i en intervju som inte kan ha undgått någon på grund av den intervjuades auktoritet , nämligen jacques delors .
vi måste därför se till att man vid regeringskonferensen verkligen diskuterar hur man skall förstärka unionens demokratiska bas , hur man skall förstärka - och det har vi redan diskuterat i denna kammare , i samband med situationen i österrike - systemet av principer , värderingar , rättigheter som ligger till grund för unionen , den roll som de politiska institutionerna skall spela inom unionen , även när det gäller att styra ekonomin .
vi litar på det portugisiska ordförandeskapet , vi litar på oss själva och vi litar på kommissionen , för allt detta kan man diskutera på ett konstruktivt och produktivt sätt under regeringskonferensen .
herr talman ! endast ett förstärkt europa kommer att klara utvidgningen .
endast ett förstärkt europa är osårbart för politiska opportunister som använder sig av ofred .
därför behövs det grundliga reformer och alltså en utvidgad dagordning för regeringskonferensen .
det finska ordförandeskapet lyssnade endast till minimalistiska regeringar och var tyvärr stendövt för det här parlamentet .
portugal kan av sina finska föregångare lära sig hur det inte skall gå till .
det är mycket viktigt att europaparlamentet och kommissionen gör gemensam sak vid den här regeringskonferensen .
de har i många fall samma intressen och samma insikter .
en väsentlig del av den gemensamma insatsen måste i alla fall vara parlamentets medbeslutanderätt vid de kommande fördragsändringarna .
av alla prioriteter så är det de som väger tyngst .
det betyder också att parlamentets ordförande och de två företrädarna måste kunna delta på en jämlik politisk nivå , alltså inte bara i arbetsgruppen utan på samma politiska nivå som kommissionen .
det finns inget som helst skäl till att folkvalda företrädare skulle delta på en lägre nivå än kommissionen .
de grundliga reformerna är vi inte bara skyldiga de nya medlemsstaterna utan även oss själva .
om vi låter europa urvattnas på grund av utvidgningen så drunknar vi i vårt eget politiska träsk .
herr talman ! det finns dagar då jag verkligen inte förstår mig på detta parlament som finner en masochistisk njutning i självstympning .
efter att på eget initiativ ha begränsat sitt deltagande i regeringskonferensen till två små platser avstår parlamentet i dag från att komplettera dagordningen för denna regeringskonferens .
oavsett om det beror på svaghet eller dumhet , och ingen av dessa möjligheter är särskilt lysande det måste ni erkänna , överger vårt parlament , genom att skynda sig att yttra sig , den enda drivkraft som fördraget ger , dvs. att kräva en fullständig dagordning för regeringskonferensen innan man uttalar sig .
varför skall vi brådskande rösta om detta yttrande i morgon den 3 februari när vi i vår styrkeposition kan vänta tills sammanträdet i strasbourg öppnas den 14 februari , och på så sätt påtvinga rådet en dagordning som äntligen är fullständig och därmed enhetlig ?
det krävs en hel del hyckleri för att dölja vår svaghet i dag .
hyckleri för att i vår resolution allvarligt beklaga att regeringskonferensens dagordning inte är i nivå med vad som står på spel , medan vi med en skyldig naivitet gör allt för att undvika att tvinga fram denna ambitiösare dagordning .
om det i slutet av denna regeringskonferens föreligger ett demokratiskt tomrum , då säger jag att de politiska grupper som velat ha denna brådska blir ansvarig för detta .
vare sig man vill det eller ej kommer besluten att förskjutas mot de femton staterna i unionen , eftersom vårt parlament självt kommer att släcka den enda strålkastare som gjorde det möjligt att något lysa upp debatterna .
jag uppmanar därför ledamöterna bland den enorma majoritet i parlamentet som i november ansåg att europas framtid förtjänade bredare debatter än reliken från amsterdam , att greppa sin vallfärdsstav och gå och övertyga sin regering om att vi måste utvidga denna regeringskonferens eftersom resolutionen från europeiska rådet i helsingfors tillåter det .
på grund av situationen i österrike är denna dag en mörk dag för europa .
man inser då att demokratins seger aldrig är vunnen och att vi måste övertyga och övertyga igen .
för att bekräfta våra grundläggande värderingar är det brådskande att skriva dem och utöver denna regeringskonferens tror jag att vi är skyldiga europa en konstitution .
herr talman ! i det förslag till resolution som vi nu diskuterar krävs precis som tidigare att den kommande regeringskonferensen skall ha en bred dagordning med genomgripande reformer av institutionerna .
som argument för detta används den kommande utvidgningen av unionen .
jag är övertygad om att det är en felsyn .
ett federalt och centralistiskt eu som styr alltmer i medlemsländerna har i själva verket sämre förutsättningar att utvidgas .
ett flexibelt eu som koncentrerar sig på färre men viktiga områden och respekterar nationella olikheter och den nationella demokratin har bättre förutsättningar att omfatta betydligt fler länder .
i resolutionsförslagets punkt d krävs en mer samordnad och öppnare ekonomisk politik på eu-nivå .
att tala om det är dock inte möjligt utan att samtidigt prata om den monetära unionen .
i den här texten sägs ingenting om de stora demokratiska och politiska problemen med valutaunionen och centralbanken - det är inte hållbart .
vill man göra eu mer demokratiskt , måste emu : s hela konstruktion omprövas .
centralbanken måste ställas under politisk kontroll , så att valutapolitikens inriktning kan styras av politiska mål som hög sysselsättning och välfärd ; insynen i centralbanken måste förbättras för att detta skall bli möjligt .
stabilitetspaktens stela och misslyckade monetarism måste omprövas och förkastas , för att vi skall kunna ha en enhetlig politik som sätter välfärdsmålen främst .
fördragets artikel 56 , som förbjuder varje ingrepp i den fria rörligheten för kapitalet , valutaspekulationen , måste tas bort så att den skadliga valutaspekulationen kan hejdas genom politisk kontroll .
i flertalet eu-länder sitter i dag regeringar som domineras av socialdemokrater .
det är anmärkningsvärt att ingen av dem kräver någon förändring i valutaunionens inriktning , nu när de har möjligheten .
det skadar ju också trovärdigheten , när man påstår att valutaunionen skulle kunna utgöra en motvikt mot det globaliserade kapitalet .
i resolutionen kräver man att europaparlamentet skall få ökat inflytande över regeringskonferensen .
det är emellertid viktigt att understryka att regeringskonferensen är och skall vara en konferens mellan medlemsstaterna .
det är medlemsländernas parlament , eller folk i folkomröstningar , som skall styra fördragets utveckling .
det är därför uteslutet att europaparlamentet ges något formellt inflytande i förhandlingsprocessen eller ratificeringen .
herr talman ! utskottet för konstitutionella frågor har föreslagit en text som i allt väsentligt är positiv , som jag kommer att rösta för , även om jag själv föreslog många ändringsförslag .
det som under alla omständigheter har hänt under senare tid visar att alla de som riktade kritik mot hur utvidgningen och revideringen av fördragen planerades hade rätt .
man kan inte utvidga unionen med 28 nya medlemmar utan att ta upp frågan om europa har några principer , några gemensamma värderingar , om europa reduceras till ett ekonomiskt frihandelsområde eller om det i stället har större ambitioner än så : att vilja vara en övernationell union , på ett sätt som måste definieras , som vill lägga ut ett nytt spår i världen mot humanitet och demokrati .
det är detta vi önskar och menar när vi kräver en europeisk konstitution .
i stället har ändringen av fördragen begränsats till en revision av vissa interna regler , en nödvändig och viktig revision , men en som inte besvarar den grundläggande fråga som ställts : vad är europa , vilka är dess gemensamma principer och därmed också dess mål och gränser ?
men politiken hämnas och även om den kastats ut från fönstret i en debatt om en begränsad dagordning , så kommer den i själva verket tillbaka genom bakdörren , och i fallet österrike genom ytterdörren , för i österrike kommer ett parti till makten som tycks verka för intolerans , främlingsfientlighet , olika former av rasism .
och det handlar inte om banden med det förflutna , detta är ett problem inför framtiden , och inget kunde vara felaktigare än att vi i den här frågan splittras mellan höger och vänster .
jag tillhör en värld , de liberala katolikernas värld , som inte hör till vänstern men som står lika fast när det gäller försvaret av värden som tolerans , de gemensamma europeiska värderingarna , som alla andra och som vägrar ha något att göra med strömningar som förnekar sådana värden .
rådet gjorde rätt som tog upp den här frågan i europa och i världen och om vi inte fäster dessa värden i ett fördrag om grundläggande rättigheter , i en europeisk konstitution , så bygger vi upp ett europa som inte har några fasta och hållbara grundvalar .
jag vet , kommissionär barnier - eller åtminstone så tror jag mig veta - att ni och samtliga företrädare för det portugisiska ordförandeskapet delar dessa värderingar : utnyttja de öppningar som kom från konferensen i december för att ta upp dessa frågor och dessa principer , för endast så kan vi konstruera ett hållbart europa .
herr talman ! jag befinner mig i den glädjande situationen att jag kan hänvisa till ett par betydelsefulla inlägg från en liten grupp av nordiska skeptiker och motståndare till den våldsamma och övergripande integrationsprocess som i grunden hotar hela det demokratiska europa .
jag tänker på inläggen från bonde och sjöstedt , i vilka de påpekar att processen innehåller en rad förhållandevis aningslösa men tveklöst rationella och maktdikterade åtgärder i riktning mot ett centralistiskt och federalt eu .
de tog helt riktigt upp problemet med den monetära unionen och den centralistiska styrningen och ställde några alternativa demokratiska principer mot denna .
jag kan tillfoga att all rationell politisk agitation i mitt hemland , danmark , går ut på att när vi utvidgar kretsen av eu-länder till detta gigantiska antal , vi utvidgar alltså bredden , så kan vi inte samtidigt integrera mer på djupet - alltså genomföra en mer intensiv kvalitativ integration mot europas förenade stater .
men det är precis det som sker .
vi har i samband med varje geografisk utvidgning av eu : s område sett att utvidgningar på bredden har följts upp av intensiva utvidgningar på djupet , och det är precis det som utskottets resolutionsförslag handlar om , särskilt punkt 7 i vilken det står att man skall ha en mer omfattande integration på djupet , och mot bakgrund av de senaste dagarnas utveckling kan man fråga sig vad vi egentligen skall ha dessa regeringskonferenser och fördragsändringar till , när regeringscheferna - i realiteten ministerrådet - fattar beslut i förhållande till en självständig medlemsstat , vilket innebär att man intervenerar i denna medlemsstats demokratiska process .
man kan tycka vad man vill om jörg haider , och personligen tycker jag att han är en mycket farlig politisk person , men man kan ju inte intervenera i ett självständigt och vänligt sinnat lands demokratiska process .
när vi genomför regeringskonferenser och bedömer om vi skall genomföra fördragsändringar , måste vi ta hänsyn till att eu utvecklas varje dag , även i strid med fördraget som vi just har sett .
jag hälsar kommissionär barnier och det portugisiska ordförandeskapet välkomna här denna eftermiddag .
den 14 februari inleds regeringskonferensen som skall avslutas i slutet av år 2000 .
detta är en stor uppgift men den kan genomföras .
jag tror att man allmänt inom alla grupper är överens om här denna eftermiddag att dagordningen i helsingfors inte kommer att räcka till för att man skall hinna med det nödvändiga reformarbetet för att förbereda europa inför utvidgningen .
med andra ord vi måste täcka mer än vad som man har kallat de viktiga &quot; amsterdamresterna &quot; .
dessa innefattar utökad användning av omröstning med kvalificerad majoritet - i mitt land godkänner vi det , men inte när det gäller beskattningsfrågor - ny röstviktning i rådet för att gynna större stater samt antalet kommissionärer i ett utvidgat europa .
vad gäller den sista punkten vill irland behålla rätten att nominera en fullvärdig och likvärdig ledamot av kommissionen utan hänsyn till det antal medlemsstater som ansluter sig .
vi är beredda att överväga en ny röstviktning i ministerrådet , under förutsättning att de större medlemsstaterna är villiga att gå med på att varje medlemsstat får en fullvärdig och likvärdig ledamot i kommissionen .
jag tror att jag talar för många mindre länder när jag hävdar den speciella åsikten .
under regeringskonferensen behöver vi även debattera om en eventuell uppdelning av fördragen i två delar - en policydel och en konstitutionell del .
vi kan godta uppdelningen av fördragen under förutsättning att det inte skulle begränsa den kontrollmöjlighet de mindre medlemsstaterna hade om omförhandlingen av fördragets alla politikområden .
med andra ord om vi inte är helt företrädda i kommissionen kommer vi inte att kunna medverka i politiska diskussioner .
således bevakar vi hela den frågan ytterst noga .
vi ser fram emot stadgan om grundläggande fri- och rättigheter och att se dess innehåll .
i amsterdamfördraget , herr talman , fastställs antalet ledamöter i europaparlamentet till 700 och en debatt behövs i detta parlament om hur det antalet skall fördelas inom ett utvidgat europa .
jag rekommenderar varmt att vi röstar igenom dimitrakopoulos och leinens resolution . i resolutionen uttrycks tydligt såväl vår besvikelse över dagordningens otillräcklighet som vår vilja att regeringskonferensen skall klaras av så snabbt som möjligt .
det framkommer för övrigt av den positiva tidtabell som vi har beslutat om .
jag anser att europaparlamentet , med de nuvarande fördragsreglerna , inte skulle ha mycket att vinna på en konfrontationspolitik .
tvärtom bör vi koncentrera oss på att utarbeta övertygande förslag för de nödvändiga reformerna , i samarbete med kommissionen , vars förslag är värdefulla .
vi måste utnyttja dialogen på alla politiska nivåer , inbegripet , naturligtvis , dialogen på de nationella parlamentens nivå .
därigenom kommer vi att skapa ett samarbetsklimat som påverkar reformens kvalitet positivt .
parlamentets företrädare på regeringskonferensen bör göra klart för förhandlingsparterna att vi framför oss , med de institutionella förändringarna för unionen , har ansvaret för unionens konstitutionella utveckling .
de måste därför inse att man inte beslutar om frågor av detta slag enbart med köpslagningslogik .
frågorna för denna regeringskonferens är väldigt känsliga .
det är möjligt att det är lätt för oss att lägga fram lösningar , frågan är dock hur bra dessa lösningar klarar av historiens granskning .
jag vill betona två punkter som kan ge upphov till spänningar .
den ena gäller den balans som fram till i dag har bevarats mellan de stora och de små staterna .
europa är inte , och kan inte heller bli , en klassisk federal stat .
de lösningar som vi väljer måste ligga i linje med europeiska unionens grundläggande logik , som är en förening av stater och den förening av folk .
det andra området där det finns risk för kollisioner är svårare .
vi kräver av den framtida europeiska unionen , på grund av den förestående ökningen av antalet medlemmar , att organen skall vara effektivare .
det betyder att de skall fungera enklare och snabbare .
europeiska unionen är dock av sin natur - och kommer så att förbli - en sammansatt och komplex flerstatlig institution .
möjligheter till påskyndande och förenkling existerar .
naturligtvis existerar de , men det finns gränser .
om dessa gränser överskrids på grund av en ensidig effektivitet , kommer europeiska unionens rättsliga grund att ha brutits ned .
jag är emellertid optimistisk .
herr talman ! regeringskonferensens mandat måste utvidgas .
den viktigaste frågan som bör läggas till är unionens interna differentiering .
det är beklagligt att man knappt ens här i europaparlamentet än så länge alls satt sig in i unionens interna differentiering som ändå är nödvändig för att unionen skall kunna utvidgas på det sätt som beslutats .
kommissionens förre ordförande jacques delors har i offentlighetens ljus på nytt lyft fram tanken om en europeisk konfederation .
han har också talat om att avant garde-länderna som ligger i täten för integrationen borde kunna gå framåt i snabbare takt än de andra och att de för klarhetens skull borde ha egna institutioner .
kommissionens nuvarande ordförande prodi och höge representanten solana har framfört liknande tankar .
europeiska liberala , demokratiska och reformistiska partiets grupp tog ställning till unionens interna differentiering genom en ståndpunkt som gruppen godkände i november i fjol och där man för europeiska unionen föreslog ett system av cirklar med en gemensam medelpunkt , &quot; en lökmodell &quot; .
i nästa resolution om regeringskonferensen måste parlamentet på allvar sätta sig in i frågan om differentiering och flexibilitet .
såväl utvidgningen som integrationens landvinningar är hotade om vi inte kan skapa ett system av cirklar med en gemensam medelpunkt .
mina kollegor frassoni och onesta har redan ganska skeptiskt tala om några aspekter av den aktuella frågan .
jag vill tillägga att jag är bekymrad över frågan om subsidiaritet , inte bara mellan union och medlemsstater utan mellan medlemsstater och deras egna internt självstyrande regioner .
denna fråga har fått otillräcklig uppmärksamhet och här finns många bekymmersamma frågor .
jag vill särskilt fästa er uppmärksamhet på en av utvidgningens följder för detta parlament .
maximalt 700 har föreskrivits som den högsta antal som detta parlament kan bestå av utan risk och för att kunna förbli en rådgivande församling .
om man tillämpar den nuvarande principen för avvikande proportionalitet , sex platser för varje stat och sedan en plats för varje halvmiljon innevånare har man redan situationen där luxemburg med 367 000 innevånare har fler ledamöter i denna kammare än wales som är en delvis självstyrande region i förenade kungariket .
skottland , med en befolkning på 5 miljoner , har åtta platser i denna kammare för ögonblicket ; danmark och finland , med samma befolkningssiffra , har sexton .
vad kommer att hända om vi bibehåller en gräns vid 700 och för in 26 procent mer befolkning med tiden och sedan antar kommissionens som jag anser dåligt övertänkta förslag att det borde bli en europeisk kandidatlista .
vad kommer att hända med ett land som skottland , som jag företräder här ?
det kommer att bli helt osynligt !
ledamöter i denna kammare bör under dessa omständigheter inte alls bli överraskade om människor i skottland och andra sådana länder vad gäller dessa diskussioner efterfrågar om utvidgning inte också borde innebära att nya medlemsstater inifrån redan existerande medlemsstater skall kunna ansluta sig .
en växande opinion i skottland är av den åsikten .
herr talman ! påståendet att europeiska unionen står i ett vägskäl innebär inget nytt .
det är ett påstående som har upprepats vid flera tillfällen .
men den här gången är det sant : vi har infört - något som är oerhört positivt - den gemensamma valutan och nu står vi inför en utvidgning .
frågan är bara : skall vi vara förberedda eller ej när vi närmar oss en utvidgning ?
är vi på väg att utvidga utan att gå grundligt tillväga eller är det just det vi gör genom att utvidga ?
det är det som är frågan och dit leder varje diskussion beträffande regeringskonferensen , dess dagordning och metoder .
det är uppenbart att rådet för ögonblicket inte har valt att utvidga genom att gå grundligt tillväga .
det innebär en fara för utvidgningen .
farligt , sett ur perspektivet av en politisk union , och givetvis svårt att förstå för allmänheten .
i rådet bör man vara medveten om att man måste gå betydligt längre på nästa regeringskonferens , om man i framtiden vill ha en väl förberedd utvidgning av europeiska unionen .
rådet rådfrågar oss och parlamentet lämnar sina synpunkter .
vi vill ha en regeringskonferens , men inte denna .
är det nödvändigt med en regeringskonferens ?
ja , naturligtvis . men inte den här typen av regeringskonferens .
man måste gå betydligt längre vad dagordningen beträffar , man måste vara betydligt djärvare i de frågor som tas upp under regeringskonferensen som måste erbjuda en ökad insyn och demokrati .
en ökad demokrati innebär att europaparlamentet i högre grad tillåts medverka , att kommissionen i större - ja i större - utsträckning får utöva sin initiativförmåga .
och givetvis att tydliga mål sätts upp .
den funktionalistiska metoden har spelat ut sin roll , på gott och ont .
så här långt har vi kommit med den funktionalistiska metoden .
har vi uppnått några resultat ?
jo då , men det gäller att ta ett kvalitativt språng , och det innebär i politiska termer , herr tjänstgörande rådsordförande , , att övertyga gemenskapens medlemmar om att det värsta vi nu kan göra är att inte uppnå målet .
herr talman , mina damer och herrar parlamentsledamöter ! på det här stadiet och efter den debatt som jag lyssnat till mycket uppmärksamt och med stort intresse , skulle jag vilja göra några kommentarer som kompletterar de riktlinjer eller anföranden som jag redan haft äran att hålla för er de senaste veckorna , vid ordförande prodis sida .
herr talman , mina damer och herrar ! era två föredragande , dimitrakopoulos och leinen , föreslog i det betänkande de lagt fram efter ett mycket exakt och seriöst arbete , att parlamentet skulle anta ett formellt yttrande enligt artikel 48 i fördraget och att regeringskonferensen med hjälp av detta yttrande effektivt kan inledas den 14 februari , såsom det portugisiska ordförandeskapet föreslagit .
i vårt ställe , och efter att utifrån samma artikel 48 i fördraget ha åstadkommit det yttrande som förväntades från kommissionen , är vi glada över att konferensen därför kan inledas , för övrigt tidigare än vad man ursprungligen tänkt .
vi vet , jag vet , att alla de veckor vi har framför oss kommer att vara nyttiga veckor .
jag skulle bara vilja göra några kommentarer efter att ha läst detta förslag till yttrande , och efter att ha lyssnat till talarna från de olika grupperna .
mina damer och herrar ! till att börja med förstår kommissionen den oro som flera av er uttryckt när det gäller omfattningen dagordningen för konferensen .
jag förstår denna oro , denna fruktan att dagordningen skall vara alltför tvingande och det förefaller mig ändå som om vi kan arbeta , såsom jag sade till utskottet för konstitutionella frågor efter helsingfors , på grundval av detta mandat från helsingfors .
det är just i den andan och inom ramen för detta mandat , men genom att använda alla fraser , allt som står skrivet mellan raderna i detta mandat , som kommissionen själv arbetat för sitt eget yttrande .
vi är inte begränsade till vad man , för övrigt oriktigt , kallar de tre resterna .
precis som richard corbett tycker jag inte heller om ordet &quot; rester &quot; , som ger en känsla av att det handlar om tre små frågor eller frågor utan betydelse .
det handlar om tre mycket allvarliga , viktiga och svåra frågor , så svåra att det kollektiva politiska modet svek oss för att behandla dem på djupet i amsterdam .
när det gäller oss - jag svarar seguro , som nyss oroade sig på den punkten - har vi inte nöjt oss med dessa tre frågor , även om jag anser att de är de viktigaste och att vi nu måste behandla dem .
de är de första , de är inte de enda frågorna , herr parlamentsledamot , som konferensen måste behandla .
vi har behandlat andra frågor och vi har tagit upp idén att andra frågor borde behandlas under denna konferens , om det portugisiska ordförandeskapet till att börja med vill , och sedan det franska , med tanke på allvaret i det vi upplever före utvidgningen .
vi är beredda att göra det , vare sig det handlar om stadgan om de grundläggande rättigheterna , där arbetet påbörjats , eller om gusp och de institutionella konsekvenserna av förhandlingarna som ägt rum om försvarspolitiken , eller om en mycket svår fråga som vi fortsätter att arbeta med , nämligen omorganisationen av fördragen .
jag har hört många kommentarer om kommissionens yttrande , som tog upp alla dessa frågor och som behandlade många av dem grundligt , inbegripet exakta demonstrationer av förslag till nya artiklar , men ingen har sagt att vi befinner oss utanför mandaten från helsingfors .
det är därför beviset på att man samtidigt som man respekterar mandatet kan , genom att använda allt det som skrivits i mandatet och alla de öppningar det innehåller , gå till botten med frågorna .
när det gäller europaparlamentets deltagande i arbetet med konferensen tror jag att minister seixas da costa är överens med mig , eftersom vi har en gemensam erfarenhet , när jag säger att det skulle vara fel av er att strunta i nivån med diskussions- och förhandlingsgruppen där era två företrädare , professor tsatsos och elmar brok , kommer att arbeta .
de sista skiljeförfarandena kommer naturligtvis , såsom alltid är fallet i varje institutionell förhandling , att äga rum och jag tror att det är bra , inom rådet och framför allt bland stats- och regeringscheferna , som kommer att ha framgången för denna konferens i sina händer .
jag vill också i förbigående påpeka att kommissionens ordförande prodi ingår i rådet och han har för avsikt att utnyttja denna plats och denna roll , vid stats- och regeringschefernas sida , bl.a. under slutperioden . men vi måste noga förbereda detta arbete i rådet .
mina damer och herrar parlamentsledamöter !
vi får alltså inte bortse från detta förberedelse- och förfiningsarbete som jag , genom min erfarenhet från amsterdam , vet är mycket viktigt och användbart , och man skall inte bara nöja sig med tekniska preciseringar .
jag tror att de personliga företrädarna för utrikesministrarna , era två företrädare och jag själv som företrädare för kommissionen , kommer att gå till botten med saken , men det blir senare , på en annan nivå , där vi också skall delta , som de sista skiljedomarna kommer att genomföras .
under hela denna konferens , mina damer och herrar , är det inte bara ställningen för förhandlarna som är viktig , utan kvaliteten i vad de säger .
och jag vill än en gång med tanke på mina erfarenheter från amsterdam inför parlamentet upprepa , oavsett vilken tvetydig eller svag ställning de två företrädarna från europaparlamentet har , att före amsterdam var kvaliteten i vad guigou och brok sade av stor betydelse i denna förhandling .
jag är säker på att det blir samma sak när det gäller mig , på min plats , och jag skall se till att idéerna från era två företrädare uppmärksammas och respekteras under hela förhandlingen .
jag är säker på att europaparlamentet då inte blir åskådare till denna förhandling , på samma sätt som kommissionen inte heller blir det .
mina damer och herrar parlamentsledamöter ! vi väntar därför med stort intresse på ert yttrande senare där ni kommer att precisera prioriteringar och konkreta förslag från parlamentet inför förhandlingen .
det är av stor vikt att de två europeiska institutioner som kommer att närvara vid dessa förhandlingar , kommissionen respektive europaparlamentet , vid sidan av rådets medlemmar , alltid och varje dag tydligt förklarar för medborgarna i unionen vilka frågor som står på spel under denna konferens och vilka svar vi förespråkar som europeiska institutioner , med ansvar för att se till att denna utvidgade union fungerar korrekt och i allas intresse .
mina damer och herrar parlamentsledamöter ! under de kommande månaderna kommer alltså kommissionen att arbeta i nära samråd , och på ett intelligent sätt , med era två företrädare , professor tsatsos och elmar brok , för att närma våra ståndpunkter till varandra , om det behövs .
sannolikt kommer våra ståndpunkter och våra positioner inte alltid att vara desamma , det kommer säkerligen att föreligga skillnader , vilket är normalt .
det som är viktigt , är att det föreligger enhetlighet , det är för att arbeta med denna enhetlighet som jag redan från början engagerat mig i mitt ämbete inom kollegiet .
vi har alltså strävan och ambitionen , i ett mycket stort antal frågor , att befinna oss på samma våglängd och höja förhandlingen .
det är ingen tillfällighet eftersom , jag upprepar det , det förefaller som om vi har samma ambition för denna förhandling och vi känner tillsammans att den verkligen utgör en sanningens minut för europeiska unionen .
herr ordförande ! jag skulle slutligen litet snabbt vilja göra tre kompletterande kommentarer .
till att börja med för att lyckönska och tacka ordförande napolitano och utskottet för konstitutionella frågor för det mycket starka och originella initiativ som togs i går genom att samla kvalificerade företrädare från de nationella parlamenten , utskottet för konstitutionella frågor och kommissionen för en första gemensam debatt .
denna dialog mellan de nationella parlamenten , europaparlamentet och oss själva är mycket viktig .
jag sade för övrigt att jag skulle ta mitt ansvar genom att själv besöka samtliga nationella parlament .
i morgon kommer jag att vara i london .
om två veckor är jag i berlin .
om tre veckor i paris , och sedan skall jag fortsätta , huvudstad för huvudstad , att i min tur delta i denna dialog .
jag finner det mycket positivt och jag ville tacka er för att ni tagit detta initiativ .
ytterligare några ord för att tacka det portugisiska ordförandeskapet och särskilt herr seixas da costa , för hans voluntarism .
det han nyss sade visar tydligt på den voluntarism och den oro som också han har : det portugisiska ordförandeskapet kan inte vara ett mellanliggande ordförandeskap .
det är detta ordförandeskap som skall inleda förhandlingen .
vi vet mycket väl att den inte kan avslutas under dessa sex månader och att det franska ordförandeskapet sedan skall ta över , med förhoppningen att det skall avsluta förhandlingen innan år 2000 är slut .
och inte bara avsluta , utan också lyckas med den , vilket inte är riktigt samma sak .
att avsluta en förhandling är inte detsamma som att lyckas med den .
ordförandeskapet kommer att ha överlämnats , men under vilka förhållanden detta överlämnande sker av er själv , herr ordförande , och av det portugisiska ordförandeskapet , blir mycket viktigt , liksom hur det sker .
det är det arbete som vi skall genomföra tillsammans , och bl.a. med impulser från er , under några månader , vilket är mycket viktigt .
vi hyser stort förtroende för er och vi har stora förväntningar på det sätt som det portugisiska ordförandeskapet , från ett litet land - men även om man är liten kan och bör man ha stora ambitioner - kommer att genomföra denna uppgift .
efter att ha lyssnat till premiärminister guterrez , utrikesministern och er själv , hyser jag detta förtroende för ambitionen hos det portugisiska ordförandeskapet och det mycket voluntaristiska sätt som det kommer att föra denna förhandling på .
ordförandeskapet kan under dessa månader räkna med kommissionens partnerskap .
slutligen , jag upprepar det , har vi en mycket stor ansträngning framför oss för att popularisera frågorna i denna förhandling .
det är svåra frågor . det är frågor om institutionell politik och mekanik som inte alltid är lätta att förklara .
det är ytterligare en anledning till att ledamöterna i europaparlamentet , ministrar och kommissionärer bör ägna litet tid åt att förklara för medborgarna och bedriva en offentlig debatt .
kommissionen kommer för sin del att ta initiativ , mina damer och herrar , till att inleda och föra denna debatt .
utförande av tjänster över gränserna
herr ordförande , herr kommissionär , värderade kolleger ! till att börja med måste jag be om ursäkt för att jag är litet hes i dag , men som österrikisk ledamot har man haft mycket att förklara och tala om i dag .
jag vill först tacka kommissionen så hjärtligt för det initiativ som den har tagit , och för de båda förslag till direktiv som vi diskuterar här i dag .
den åtgärdar därmed två graverande brister på den inre marknaden som är av stor betydelse för det europeiska näringslivet och för 5 miljoner tredjelandsmedborgare i europeiska unionen , vilka är här som arbetstagare eller som individer .
dagens situation , och det bör man än en gång betänka , ser ut så att det i fråga om arbetstagarna visserligen föreligger domar från eg-domstolen , i synnerhet domen som gäller rush portuguesa och van der elst .
de har visserligen klarlagt att friheten att tillhandahålla tjänster måste medge att man använder sig av tredjelandsmedborgare som arbetstagare för gränsöverskridande tjänster , och detta även utan att kunna utverka arbetstillstånd .
frågan om viserings- och uppehållsvillkor fördes inte utförligen på tal , och inte heller medlemsstaterna kunde sedan förklara denna fråga .
men inte heller med hänsyn till bortfallet av arbetstillståndet har alla medlemsstater hållit sig till domstolens domslut utan upprätthåller fortfarande i dag en mängd otillåtna barriärer för gränsöverskridande tjänster , barriärer som ofta är omöjliga att övervinna , i synnerhet för små företag .
för de egna företagarna ser situationen så ut att gemenskapens nuvarande regelverk inte föreskriver någon rätt för tredjelandsmedborgare att utföra gränsöverskridande tjänster .
här behöver man i varje fall en rättsakt .
båda förslagen till direktiv syftar till att underlätta friheten att tillhandahålla tjänster för eu-företag .
det handlar inte om nya rättigheter för tredjelandsmedborgare , som efterbildar den fria rörligheten .
alla bestämmelser , inresa och frågor som gäller uppehållet , skall betraktas som tillägg till denna frihet att tillhandahålla tjänster .
tillsammans med utskottet för rättsliga frågor och den inre marknaden anser jag därför att den av kommissionen valda rättsliga grunden är riktig och att den motsatta åsikt som företräds i utlåtandet från rådets rättstjänst inte är tillämplig .
jag ser därför inte heller något verkligt hinder för att båda förslagen till direktiv snabbt skall kunna vidarebehandlas i rådet .
jag tror också att de av parlamentet föreslagna ändringarna bör göra att direktiven lättare blir antagna i rådet , jämfört med kommissionens förslag .
många av våra ändringar går tillbaka till betänkligheter som även yttrats i rådet , och vi försöker att förena dessa betänkligheter med det uppdrag som gällande rätt och ekonomiskt förnuft ger oss .
även med tanke på acceptansen i rådet kan jag bara vädja till kommissionen att så snart som möjligt fullständigt överta de ändringar som parlamentet antagit , även om de delvis avviker avsevärt från kommissionens ursprungliga förslag .
jag är fast övertygad om att vi på denna grundval lättare kan uppnå enighet i rådet .
nu till de viktigaste ändringarna som vi föreslår . en väsentlig skillnad består i att vi i stället för ett system med frihet att tillhandahålla tjänster plus anmälning av varje enskilt uppdrag inte längre räknar med möjligheten att man för varje enskilt uppdrag skall kunna begära att det i förväg anmäls till det mottagande landet .
detta system förefaller oss oanvändbart i praktiken .
som kompensation för detta måste dock , innan eg-kortet för tillhandahållande av tjänster ställs ut , alla eventuella hinder ha undanröjts , och gentemot kommissionens förslag måste skärpta villkor ha uppfyllts för att eg-kortet för att tillhandahålla tjänster skall kunna ställas ut .
kraven på vederbörlig sysselsättning , legalt uppehåll och försäkringsskydd måste finnas inte bara vid tidpunkten då eg-kortet ställs ut , utan under hela kortets giltighetstid , plus tre månader därefter .
därigenom bör den mottagande staten ha en garanti för att arbetstagaren respektive den egna företagaren efter fullgjort uppdrag också återvänder till den stat han kommer från , och i händelse av sjukdom och olycksfall täcks av försäkringar .
inresan och situationen som rör uppehållstillståndet skall också ha klarlagts innan kortet för tillhandahållande av tjänster ställs ut , nämligen inom ramen för ett överklagandeförfarande .
vi föreskriver att eg-kortet för tillhandahållande av tjänster inte måste begäras för alla medlemsstater , utan att det också kan begäras för enskilda medlemsstater .
jag tror att detta system också bättre motsvarar de praktiska behoven .
samma sak hoppas jag man åstadkommer genom förslaget att sänka minimilängden för den tidigare sysselsättningen till tre månader , och att inrikta giltighetstiden för kortet för tillhandahållande av tjänster beroende på längden på den tidigare sysselsättningen på ett flexibelt sätt .
men vi anser fortfarande att den maximala giltigheten för kortet för tillhandahållande av tjänster skall ligga vid 12 månader .
vad gäller de egna företagarna föreslår vi också , som tillägg till de redan beskrivna ändringarna , att etableringskriteriet måste skärpas och att vi föreskriver en möjlighet att bemöta ett eventuellt missbruk på grund av falskt egenföretagande .
jag vill också kort gå in på föreliggande ändringsförslag , som går utöver ändringsförslagen från utskottet för rättsliga frågor och den inre marknaden .
jag vill naturligtvis också säga att jag även i fortsättningen stöder de av detta utskott framlagda ändringarna , som antogs enhälligt i utskottet .
jag har själv för min grupp lämnat in fyra ändringsförslag , som väsentligen hänför sig till det korrekta sättet att citera ett beslut från rådet .
jag måste säga att jag här från parlamentets tjänsteenheter har fått ytterst motsägande uppgifter om hur nu detta beslut från rådet skall citeras korrekt ; endast med nummer , endast med datum , med båda , hur utförligt det skall citeras från rådets beslut .
två ändringsförslag togs bort av tjänsteenheterna , eftersom man enligt uppgift redan tagit hänsyn till innehållit i dem i betänkandet .
jag drar tillbaka de två ytterligare ändringsförslagen - det är ändringsförslag 18 i betänkandet om egenföretagarna och 21 om de anställda .
jag kan bara vädja till talmanskonferensen att så snart som möjligt enas om hur man i fråga om kommittésystemet skall agera korrekt när det gäller citat .
det skulle underlätta livet för föredragandena i denna kammare väsentligt i framtiden .
det föreligger också ett ändringsförslag till båda betänkandena från kollegan de palacio .
jag måste tyvärr säga att jag inte kan stödja detta ändringsförslag , eftersom det skulle förändra substansen i de resultat som vi enhälligt uppnådde i utskottet för rättsliga frågor och den inre marknaden , och jag vill bibehålla det som vi i detta utskott efter långa diskussioner gemensamt kom fram till .
avslutningsvis vill jag tacka alla kolleger som har bistått mig i utskottet för rättsliga frågor och den inre marknaden i dessa inte direkt lätta betänkanden .
i synnerhet vill jag nämna kollegan wieland , som har den otacksamma rollen som medföredragande och långt utöver det vanliga tagit del i utformningen av detta betänkande med mycket bra och konstruktiva idéer , utan att få någon del av föredragandens lagerkrans .
därför vill jag här särskilt nämna det !
( nl ) herr talman ! jag är glad att jag får tillfälle att efter anförandet av föredraganden , berger , göra några inledande kommentarer varefter jag naturligtvis med allt det intresse som krävs skall lyssna till de följande talarna .
om ni tillåter , herr talman , skulle jag sedan i slutet av debatten vilja ta upp de olika ändringsförslagen mer ingående .
jag vill tala om att kommissionen gläder sig åt europaparlamentets stöd för de två förslag för tillhandahållande av tjänster och arbetstagare från tredje land , vilka debatten nu gäller .
jag är särskilt tacksam för det arbete som berger lagt ner vid behandlingen av de här förslagen som ju är politiskt känsliga och som är en politisk utmaning .
jag vill också tacka palacio så mycket för hennes mycket viktiga bidrag som ordförande för utskottet för rättsliga frågor och den inre marknaden .
kommissionen gläder sig särskilt åt parlamentets förslag om ett effektivare förfarande för utfärdande av kortet för tillhandahållande av tjänster .
när det finns möjlighet att ansöka om ett sådant kort för en eller flera eller för alla medlemsstater så blir förfarandet ännu flexiblare .
kommissionen går också med på den föreslagna giltighetstiden för kortet .
jag anser emellertid att en arbetsperiod på tre månader inte räcker som bevis för att en arbetstagare är etablerad i en medlemsstat .
kommissionen kan också gå med på en bestämmelse för de fall då arbetskontraktet mellan tjänsteleverantören och arbetstagaren plötsligt upphävs .
ett effektivt förfarande för utfärdande av kortet innebär att företag som tillhandahåller gränsöverskridande tjänster också verkligen kan utöva sina rättigheter på grund av den inre marknaden .
vi tycker att det verkar överdrivet om andra medlemsstater får möjlighet att för utfärdandet av ett kort genomföra systematiska kontroller med avseende på den allmänna ordningen .
en medborgare från ett tredje land med en legal ställning måste ju också få komma in i andra medlemsstater .
det hindrar inte dessa medlemsstater från att inom ramen för den föreslagna meddelandeskyldigheten vidta åtgärder med avseende på den allmänna ordningen .
förslaget om att uppehållstillståndet i en medlemsstat borde vara tre månader efter kortets giltighetstid kan kommissionen inte heller godta .
det är inte godtagbart att den berörda medborgaren från ett tredje land stannar längre i medlemsstaten efter det att tjänsterna tillhandahållits .
därför stöder kommissionen i båda fallen ändringsförslag 22 av palacio .
när det gäller det andra förslaget så inser kommissionen att det måste vara tydligt vad som menas med en egenföretagare och skall därför komma med en lösning i det ändrade förslaget .
det var några inledande kommentarer om de viktigaste ändringsförslagen .
jag hoppas att jag i slutet av den här debatten , när alla talare sagt sitt , får ytterligare tillfälle att ta upp de olika ändringsförslagen .
herr talman , mina damer och herrar ! ppe-gruppen kommer med stor majoritet att rösta för ändringsförslagen från utskottet för rättsliga frågor och den inre marknaden och även den ändrade versionen under morgondagen .
jag vill i mina utlägg inskränka mig till två betänkanden .
det ena gäller frågan om vad detta direktiv över huvud taget skall verka för - verka för i dess egentliga betydelse .
vi har för det första näringslivets och även de enskildas intressen .
i mina inlägg utgår jag till att börja med från att det handlar om en rättskaffens och rejält arbetande enskild .
för det andra har vi medlemsstaternas intressen , som med tanke på dem som berörs kanske också måste utgå från att det föreligger ett worst case .
om vi tänker på den ena ytterligheten , medlemsstaternas intressen , så finns det säkert goda anledningar att sätta hindren för detta eg-kort relativt högt .
sedan finns det anledning att trots detta eg-kort på ett tidigt stadium införa anmälningsplikt .
om jag tänker på den andra ytterligheten , alltså så få hinder som möjligt , då riskerar jag att jag i fråga om detta förfarande över huvud taget inte kommer att få uppleva någon lagstiftning , eftersom medlemsstaterna då inte kommer att godkänna direktivet .
resultatet blir alltså antingen att jag visserligen har ett direktiv för eg-kortet för tillhandahållande av tjänster , men , eftersom hindren för näringslivet är mycket höga , i själva verket inte har något eg-kort för någon .
i det andra fallet har jag inte alls något direktiv .
ingetdera resultatet är tillfredsställande .
kanske är detta också anledningen till , som man hör sägas , att förhandlingarna har hakat upp sig även i rådet .
nu har vi försökt att åstadkomma ett mellanting mellan det ena intresset - ordre public - och det andra intresset , och att finna en så lätt lösning som möjligt .
vi vill ha en lösning där vissa hinder för näringslivet byggs upp , men där man sedan , när dessa hinder övervunnits , uppnår en så smidig hantering som möjligt .
vi vill därför att eg-kortet för tillhandahållande av tjänster begärs för en eller flera medlemsstater .
om ett företag i frankrike säger att man har en medarbetare som ständigt måste arbeta i danmark och bara i danmark , då skall detta eg-kort för tillhandahållande av tjänster också bara begäras för danmark .
då kommer de byråkratiska hindren för detta att vara lägre .
som en motåtgärd vill vi dock att det inte längre skall finnas några fler tidiga anmälningsplikter , utan att arbetstagaren enbart skall ha med sig anledningen till arbetena i den andra medlemsstaten , till exempel i form av det avtal som ligger till grund för dem .
därför måste jag också säga att jag till slut uttalar mig för ändringsförslagen från utskottet för rättsliga frågor .
kanske finns det också hos kommissionen fortfarande kvar en viss rest av missuppfattning .
vi vill att man uppnår en helt flexibel lösning .
om en medlemsstat förklarar att man plötsligt har problem , eftersom personen har begått en stöld , man har problem , och detta eg-kort för tillhandahållande av tjänster är utställt för ens land , då kan det enskilda landet av de anledningar som finns i detta direktiv i viss mån dra tillbaka giltigheten för eg-kort , på ett flexibelt och intelligent sätt .
låt mig också helt kort gå in på en annan sak .
de flesta som hittills befattat sig med direktivet är jurister .
vi vet alla att det fortfarande finns olika beståndsdelar i fördraget , delvis mycket gamla beståndsdelar i fördraget , som fortfarande heter eg .
vi vet att detta direktiv baserar sig på eg-rätt och inte på eu-rätt .
men före valet verkade vi - rådet , kommissionen , parlamentet , pressen , fackföreningarna , organisationerna - för att detta europa skall bli mer förståeligt för medborgaren .
vi har ansträngt medborgarna genom att ändra eeg till eg till eu .
nu har man förstått eu .
vi gör oss själva och medborgaren en otjänst om vi nu döper den produkt som vi ger ut till eg-kort för tillhandahållande av tjänster och inte till eu-kort för tillhandahållande av tjänster .
för medborgaren är eu-världen intressant , det är den som gäller för honom .
jag ber rådet och kommissionen att gå i den riktningen .
herr talman ! det har blivit senare än någon av oss trodde det skulle bli när vi planerade denna session så jag skall verkligen fatta mig kort .
en av orsakerna till varför vi är försenade är för att vi använde tiden tidigare i dag till att rätteligen framföra det fast förankrade motståndet i detta parlament mot varje form av främlingsfientlighet och rasism .
detta direktiv handlar naturligtvis inte i sig självt direkt om det .
det handlar om att se till den inre marknadens behov , att skapa flexibilitet och att agera på ett förnuftigt och flexibelt sätt för att skapa sysselsättning för människor från tredje land både som anställda och som egenföretagare .
det handlar i sig själv också om att undvika att vara obefogat restriktiv mot främlingar bara för att han eller hon är en främling .
vi välkomnar det och då vi anser att det är en förnuftig och riktig bestämmelse kommer vi att stödja den mest generösa versionen som vi anser är i överensstämmelse med lagstiftningen .
( es ) - herr talman , herr kommissionär ! jag vill börja med att poängtera det utmärkta arbete som berger har gjort och även rent allmänt utskottet för rättsliga frågor och den inre marknaden , som har infört nyskapande idéer i detta direktiv som jag hoppas kommer att godkännas av kommissionen och rådet .
jag har emellertid lagt fram ett ändringsförslag .
fru berger , i ert ändringsförslag 2 , skäl 6 , tar ni upp rättssäkerheten .
den första punkt där vi har en avvikande mening är uppehållstillståndets förlängning med tre månader , för det skapar endast rättsosäkerhet .
ni har - av naturliga skäl - uttryckt er oro , som bekräftats av wieland , för möjligheten att en arbetstagare försvinner när dennes arbetstillstånd har löpt ut , men jag anser att ni samtidigt underlättar denna möjlighet i och med förlängningen med tre månader .
om giltigheten för eg-kortet för tillhandahållande av tjänster upphör ett visst datum , bör den också upphöra det datumet .
det är en förutsättning för rättssäkerheten .
å andra sidan , vad beträffar punkt d ) i ändringsförslag 10 som åsyftar det första direktivet , nämner ni att en medlemsstat på grund av allmänhetens säkerhet eller bestämmelser om den allmänna ordningen , kan vägra erkänna kortets giltighet .
redan nu sker kontroller som ex ante fastställs i artikel 4 i direktivet .
det saknar betydelse för en arbetstagare inom schengenområdet , för denne har redan genomgått en kontroll för att få resa in i den första medlemsstaten , och den andra medlemsstaten kan ex ante , om vissa skäl föreligger , neka denna arbetstagare inresa i landet .
det finns därför ingen anledning att bevara denna rättsosäkerhet .
om det inte rör sig om en schengenstat så förutses den möjligheten i sista stycket i mitt ändringsförslag 22 , i alla avseenden och med det jag anser vara en bättre rättssäkerhet .
staternas fria val som ni föreslår i punkt e ) i ert ändringsförslag 10 rimmar inte med texten i övrigt i ert utmärkta betänkande .
därför uppmanar jag er kolleger att ta del av mitt ändringsförslag , och hoppas att vi i morgon kan komma fram till en lösning .
av allt att döma tycks dessa två förslag införa vissa ändringar i förfarandena för att underlätta fri rörlighet i hela europa och för att låta de nya domstolsfall som berger refererade till i sitt öppningsanförande få effekt .
i fråga om förenade kungariket tror vi emellertid att man där går längre än så på ett sätt som är oacceptabelt .
delvis finns verklig substans delvis är det med hänsyn till den rättsliga grunden vad gäller förenade kungarikets särskilda ställning .
enligt de protokoll som finns i fördragen behåller förenade kungariket sin egen gränskontroll .
enligt det system som föreslagits på dessa lagstiftningsområden kommer medborgare i tredje land som vill flytta till förenade kungariket att enligt de beskrivna förfarandena kunna göra detta med hjälp av ett servicekort utfärdat av en annan medlemsstat och därigenom kringgå landets gränskontroller .
om det nuvarande gränskontrollsystemet i förenade kungariket skall ändras bör den ändringen göras av förenade kungarikets regering och parlament och inte i förbifarten genom det europeiska lagstiftningsförfarandet .
av det skälet skall vi rösta mot båda dessa förslag .
herr ordförande , herr kommissionär , mina damer och herrar ! först vill jag tacka föredraganden och kollegan wieland så hjärtligt för deras ansträngningar att så homogent sammanfatta de olika ändringsförslagen och de olika intressena i detta betänkande .
dessa båda förslag bidrar till att genomföra en av de fyra kärnprinciperna för den inre marknaden , fri rörlighet för tjänster .
de nya bestämmelserna för gränsöverskridande tjänster kommer utan tvivel att förbättra både den inre marknadens funktion och företagens konkurrens- och handlingskraft .
de strikta ramvillkoren för utställandet av - och här citerar jag kollegan wieland - eu-kortet för tillhandahållande av tjänster är oundgängliga , eftersom de tjänar till att förhindra missbruk , exempelvis illegal invandring och falska kontrakt .
varför anser jag att direktivet är så nödvändigt ?
av tre anledningar : på grund av den ekonomiska betydelse som arbetskraften från tredje land har i eu , på grund av företagens konkurrenskraft och på grund av den inre marknadens friktionsfria funktion .
därför välkomnar jag å ena sidan den strikta ramen , och vädjar å andra sidan om att de lämpliga kontrollerna som medlemsstaterna genomför blir så effektiva och enkla som möjligt .
min sista fråga , eftersom man alltid frågar mig om det , går till kommissionen : kommer direktivet att bli prejudicerande för anslutningsförhandlingarna ?
hur kommer artikel 1 ur er synpunkt att tolkas , eftersom detta spelar en viktig roll i anslutningsförhandlingarna och just för vårt land som gränsar till många nya länder ?
de företagare som hittills tvingades konstatera att två av de viktiga friheterna , nämligen fri rörlighet för personer och tjänster , inte gällde för dem var dock tvungna att gå igenom en oändlig byråkratisk immigrationsprocess i medlemsstater där en tjänst skulle tillhandahållas .
det finns cirka tretton miljoner medborgare från tredje land som uppehåller sig i europa .
jag utgår från att , även om det inte är känt exakt hur många av dem som är företagare , deras antal säkert inte är litet .
hittills har deras tillträde till hela europeiska unionen inte reglerats genom gemenskapsrätten .
syftet med de två aktuella förlagen till direktiv är att främja den fria rörligheten för tjänster på den inre marknaden genom införande av eu-kortet för tillhandahållande av tjänster .
jag tycker det är viktigt att i det sammanhanget understryka att utfärdandet av ett sådant kort skall ske på ett flexibelt sätt , nämligen inom fem dagar efter att en enkel förklaring lämnats till den medlemsstat där tjänsten skall tillhandahållas och att , för att undvika missbruk , den här handlingen skall ha en begränsad giltighet och inte automatiskt kunna förlängas .
jag har också med intresse tagit del av de invändningar som kommissionären fört fram här .
efter att ha studerat de inlämnade ändringsförslagen har jag också konstaterat att vi i stor utsträckning kan godta dessa invändningar och därför skall anpassa hur vi röstar efter detta vid omröstningen i morgon .
avslutningsvis skulle jag vilja tacka föredraganden berger för den noggrannhet med vilken hon undersökt de olika ändringsförslagen och på det sättet givit sitt betänkande ett viktigt innehåll .
jag tror att vi med det här betänkandet tagit ett nytt steg mot förverkligandet av den inre marknaden .
tack för att jag nu får tillfälle att mer specifikt gå in på de olika ändringsförslagen och i det sammanhanget skulle jag också vilja säga något till lord inglewood om den anmärkning han nyss gjorde .
när det gäller det första förslaget om arbetstagare från tredje länder så är kommissionen beredd att anta ändringsförslagen 2 , 11 , 12 , 15 , 16 och 22 .
även ändringsförslagen 7 och 8 är godtagbara om utstationeringssituationen i ursprungslandet kan fastställas .
kommissionen godtar också ändringsförslag 11 , förutom med avseende på den föreslagna perioden för tidigare anställning på endast tre månader . det har jag redan förklarat tidigare .
även ändringsförslag 13 är välkommet om det härigenom införs ett flexibelt tillämpningsområde för kortet från en medlemsstat till alla medlemsstater .
vad kommittésystemet beträffar så kan ändringsförslagen 14 och 21 också delvis godtas när det gäller parlamentets rättigheter .
ändringsförslag 10 kan kommissionen , tyvärr , inte godta när det gäller tremånadersperioden och den mottagande medlemsstatens roll .
kommissionen stöder i det avseendet ändringsförslag 22 , vilket jag redan påpekat .
personligen känner jag sympati för namnet &quot; eu-kort för tillhandahållande av tjänster &quot; som föreslås i ändringsförslag 1 men amsterdamfördraget tillåter inte det .
i ändringsförslag 18 hänvisas till direktiv 96 / 71 angående minimilöner som redan tillämpas , så det behövs ingen ändring .
om kommissionen skulle godta ändringsförslag 17 så skulle det innebära att en enkel anmälningsplikt skulle gälla om inget giltigt kort lämnats .
det är väl ändå i strid med intressena i samband med den allmänna ordningen i medlemsstaterna .
ändringsförslag 19 är också oacceptabelt med hänsyn till mina beaktanden kring ändringsförslag 10 .
kommissionen har samma ståndpunkt när det gäller liknande ändringsförslag till det andra förslaget .
jag vill tillfoga att ändringsförslag 10 är helt godtagbart när det gäller det förslaget .
med avseende på ändringsförslag 15 om definitionen av begreppet &quot; egenföretagare &quot; skall kommissionen , som jag redan sagt , se till att ta fram en nöjaktig lösning för att tillmötesgå de invändningar som rests .
då övergår jag till lord inglewoods anmärkning .
han hänvisade till de gränskontroller som finns med avseende på förenade kungariket och jag skulle vilja säga att ingen medlemsstat , och alltså inte heller förenade kungariket , har skyldighet att avskaffa kontrollerna vid de gränser som fortfarande finns .
det gäller , som sagt , även för belgien där den aspekten nyligen var aktuell .
angående karas anmärkning skulle jag vilja säga att jag fick intrycket att han talade om möjligheten att arbetstagare från polen utnyttjas i hans land .
kommissionen skulle vilja föreslå en lösning på det problemet varvid den lösningen skulle gälla för alla företag i europeiska unionen som anställer personal från länder utanför eu .
frågan är sedan om de två fallen skall behandlas lika .
det är en fråga som jag tycker hör hemma i debatten om europeiska unionens utvidgning och kanske inte i den här debatten .
för kommissionens räkning ställer jag mig gärna till karas förfogande om han skulle vilja ha ytterligare information i denna mycket viktiga fråga .
jag står alltså till förfogande .
avslutningsvis skulle jag vilja tacka parlamentet för den mycket konstruktiva debatten om de viktigaste aspekterna av de här förslagen och speciellt naturligtvis den viktigaste föredraganden , berger .
tack så mycket , kommissionär bolkestein .
förstainstansrätten
herr talman ! jag vill börja med att gratulera föredraganden till ett betänkande , som vid en första genomläsning endast ger intryck av att bekräfta och acceptera .
bakom det här betänkandet döljer sig emellertid ett omfattande och effektivt arbete som redan har lett till vissa resultat : handlingens införlivande i det finska ordförandeskapets löfte den 7 december 1999 om att utvidga dagordningen för regeringskonferensen till att omfatta en undersökning av de framtida förändringarna av gemenskapens domstolars organisation , sammansättning och behörighet .
därför vill jag framföra mitt erkännande av vice ordförande marinhos insats .
herr talman , en reform av gemenskapens rättsväsende har blivit en nödvändighet om man i framtiden skall kunna skipa rättvisa inom rimliga tidsramar , om europeiska unionen i framtiden vill ha en rättskipning på samma nivå som det politiska projekt som vi har påbörjat .
i dag - och det säger jag med stolthet och glädje - har vi här i parlamentet haft ett ypperligt tillfälle att visa i vilken utsträckning vi européer anser att det politiska projektet är betydligt mer än den inre marknaden , ett projekt som i större utsträckning baserar sig på principer än på ekonomiska intressen .
för bakom principerna , herr talman , döljer sig alltid rättvisan .
men justice delayed is justice denied ( att skjuta upp rättvisan är det samma som att neka den ) , och det är något vi bör fundera över .
oroväckande uppgifter framkommer av det arbetsdokument som domstolen själv har förberett .
mot bakgrund av detta är reformprojektet under föredragande av vice ordförande marinho välkommet .
denna lösning är ett lappverk , men även ett lappverk får duga , för vi kan för närvarande inte - något som han har påpekat - förvänta oss en stor reform av systemet på regeringskonferensen .
vi måste komma med lösningar som , även om de är provisoriska , bidrar till en snabbare och effektivare rättskipning .
det är två saker jag vill ta upp i det här inlägget , och som faller utanför själva betänkandet , på grund av den skyldighet som parlamentet enligt fördraget har att utarbeta ett kort och koncist betänkande utan någon fördjupning .
det är två förslag från vice ordförande marinho som , det vågar jag nog påstå , stöds av hela utskottet för rättsliga frågor och den inre marknaden .
det första innebär att domarna i förstainstansrätten skall förses med ytterligare en référendaire .
det andra är att översättningstjänsten vid förstainstansrätten skall skiljas från den vid domstolen .
i dagsläget måste förstainstansrätten vänta mycket länge på att få sina domar översatta .
vi utgör en gemenskap , vars grundläggande princip enligt fördraget är en kulturell och språklig mångfald , och vi får under inga omständigheter överväga att avskaffa en sådan viktig möjlighet som att få ta del av en dom på det egna språket .
när vi ändå talar om regeringskonferensen , låt oss då tänka på två saker .
det första gäller detta parlament .
jag tror inte det skadar att vi insisterar på en större medverkan vad domstolen beträffar , och då även i utnämnandet av domarna .
vi vill framför allt och i första hand att domstolens behörighet skall utvidgas samtidigt som förmågan att uppfylla sina skyldigheter , det vill säga dess resurser .
vi vill att behörigheten skall utvidgas , i synnerhet vad gäller avdelning iv i eg-fördraget och avdelning vi i eu-fördraget , och att man i förbifarten undersöker vissa alternativ på dessa områden som är så utomordentligt viktiga för våra medborgare .
då syftar jag åter igen på de uttalanden som vi har fått ta del av de senaste dagarna .
herr talman ! jag vill gratulera föredraganden och välkomna innehållet i detta betänkande .
det har fått mig att tänka på två problem som jag har fått nyligen i mitt eget valdistrikt .
båda gäller nära förestående avgörande i eg-domstolen .
det första fallet gäller en stor hängbro och om brotullarna för den skall vara momspliktiga eller inte .
beslutet skulle få enorma följder för vår lokala ekonomi .
det andra fallet gäller en dam som skall pensioneras inom tretton veckor och som förtvivlat väntar på ett domstolsavgörande som allvarligt kommer att påverka hennes ekonomiska villkor som pensionär .
detta är bara två exempel på verkliga vardagliga problem som förseningar i europas rättssystem skapar .
dessa förseningar kan innebära personliga svårigheter och även tragedier .
med detta säger jag inte att alla våra egna nationella rättssystem fungerar perfekt men alltför ofta kan det hända att de väntar på ett förhandsavgörande från eg-domstolen .
statistiken visar en oroande stigande trend i fråga om den tid som krävs för att hantera förhandsavgöranden .
detta skall inte ses som kritik av domstolen eller dess personal utan snarare domstolens struktur och dess brist på resurser i en växande europeisk union .
förslagen i detta betänkande är mycket välkomna som ett tillfälligt avhjälpande åtgärd , men europa är en rättslig konstruktion och dess domstolar är avgörande för att allt skall fungera på vederbörligt sätt .
i avvaktan på den kommande utvidgningen måste regeringskonferensen ta itu med grundläggande reformer och omstrukturering av domstolssystemet .
i annat fall kommer vi alla , som valda representanter , att få ta emot mer och mer högljudda krav från våra medborgare då de inte får tillgång till snabba och effektiva rättssystem .
herr talman , mina damer och herrar , kolleger ! jag vill också tacka föredraganden för detta utmärkta betänkande .
jag är också helt införstådd med hans slutsatser , där han särskilt föreslår att antalet rättssekreterare för domarna vid förstainstansrätten skall ökas och att förstainstansrätten skall ges en egen översättningstjänst .
jag anser att detta faktiskt är nödvändigt , eftersom vi vid utskottets för rättsliga frågor besök i luxemburg fick höra att , eg-domstolen , naturligtvis med naturnödvändighet , så att säga ofrånkomligt , har företräde framför förstainstansrätten vid utnyttjandet av den gemensamma översättningstjänsten , och att därför viktiga saker ofta inte kan behandlas tillräckligt vid förstainstansrätten .
men jag anser också att reformerna måste gå längre än vad vi nu kommer att besluta om .
jag tror att det exempelvis är värt att överväga att man på de områden , där redan domarkollegier , som liknar domstolar , i förväg fäller ett avgörande - jag vill bara nämna alicante eller hur nu detta har planerats för den europeiska ämbetsmannalagen - i förekommande fall gör förstainstansrätten till sista instans , och här upprättar en avslutande behörighet .
jag inser också att vi förmodligen måste göra något i samband med kommissionens tendenser att åternationalisera konkurrensavgöranden och lägga tillbaka dem på den nationella nivån .
här förefaller det nödvändigt att överväga detta , eftersom dessa fall ju då inte längre skulle hamna hos förstainstansrätten , utan som förlagor till beslut vid eg-domstolen .
vi bör överväga hur vi skall hantera denna situation .
eventuellt bör det också finnas möjlighet att lämna förlagor till beslut i konkurrensärenden till den specialiserade avdelningen vid förstainstansrätten .
dessutom måste man också överväga , om det är rätt - och vi har just haft fall , där ledamöter eller grupper har överklagat mot europaparlamentet - att förstainstansrätten är ansvarig för sådana frågor , även om det egentligen handlar om författningsfrågor och dessa saker helt logiskt egentligt hör hemma hos eg-domstolen och mindre hos förstainstansrätten .
en sista punkt : jag tror också att det behövs en demokratisk kontroll av olaf .
för ögonblicket befinner sig olaf i ett vakuum och kan göra vad den vill .
jag anser att det är nödvändigt att olaf kontrolleras av en domstol .
den enda domstol som kan göra det på ett förnuftigt sätt skulle vara förstainstansrätten .
också detta skulle vara en impuls för den fortsatta reformprocessen .
herr talman ! jag skulle vilja börja med att instämma med dem som gratulerade föredraganden för detta dokument .
europeiska unionen är ett system grundat på lagar .
den måste därför ha ett domstolsväsen för att genomdriva dessa lagar .
om domstolarna dessutom inte kan klara av den arbetsmängd som läggs på dem på ett riktigt och snabbt sätt händer det som palacio vallelersundi redan påpekat , nämligen att försenad rättskipning blir samma som nekad rättskipning .
domstolens bevis är att det händer nu och det pekar mot åtgärder som kan vidtas nu för att lindra problemet .
men som marinho påpekade , mer krävs , men det får vänta till regeringskonferensen .
i mitt eget land talas det mytiskt om de myllrande horderna av anonyma brysselbyråkrater men man talar aldrig om antalet europeiska domare .
det finns mindre än tre dussin i toppen på det europeiska rättskipningssystemet - knappast en överbemanning med tanke på deras ansvarsfulla uppgifter i hjärtat av det europeiska rättssystemet .
hur stor deras betydelse är kan man se i de politiska följderna av förseningen med att lösa den mycket viktiga engelsk-franska tvisten om brittiskt nötkött som har skapat så mycket ilska i mitt land och sådan besvikelse över unionens handläggning av domstolstvister .
detta har förvärrats , något som några av mina rådgivare anser , av procedurreglerna i de franska domstolarna som gör det nästan omöjligt för icke franska medborgare att öppna process mot den franska regeringen .
det uppfattas faktiskt som omöjligt .
detta kontrasterar mycket ofördelaktigt mot förenade kungarikets domstolar där spanska fiskare framgångsrikt lyckades väcka åtal mot förenade kungarikets regering under mycket jämförbara förhållanden .
vad som händer i frankrike , herr talman , verkar vid första anblicken vara ett fall av diskriminering mot övriga eu-medborgare på grund av nationalitet och därmed bryta mot fördragen .
jag skulle därför vilja be kommissionären , som var vänlig nog att kommentera mina inlägg i den tidigare debatten , att undersöka detta och meddela resultaten till parlamentet och mig .
jag skulle vara tacksam om kommissionären i sin slutkommentar kan bekräfta att han kommer att göra detta .
( nl ) herr talman ! å kommissionsordförande prodis vägnar skulle jag gärna vilja svara så här .
kommissionen noterar den ståndpunkt som europaparlamentet i dag intagit angående domstolens och förstainstansrättens begäran om att å ena sidan till förstainstansrätten överlåta den bedömning av vissa överklaganden som domstolen nu har ensam behörighet för och å andra sidan öka antalet ledamöter i förstainstansrätten .
jag skulle vilja tillfoga att jag för kommissionens räkning med stort intresse lyssnat till de anföranden som hållits här alldeles nyss och att jag mycket väl begriper den oro som ligger till grund för dessa anföranden .
den oron är berättigad .
det har flera gånger sagts att justice delayed is justice denied .
kommissionen begriper den inställningen .
mot bakgrund av den insikten skulle jag vilja fortsätta mitt svar på följande sätt .
som parlamentet vet så är kommissionen övertygad om att gemenskapens rättsinstanser utan en grundlig reform löper risken att på kort sikt inte längre kunna utföra sina uppdrag inom rimliga tidsfrister .
kommissionen har därför också rådfrågat en expertgrupp om de reformer som skulle kunna genomföras för att domstolen och förstainstansrätten skall behålla kvaliteten och koherensen i sina domslut under kommande decennier .
kommissionen känner till förstainstansrättens begäran om personalförstärkning men för ögonblicket anser kommissionen att den föreslagna överföringen av behörigheter skall betraktas i ljuset av den undersökning som jag nyss nämnde och kommissionen skall lämna sitt yttrande om domstolens och förstainstansrättens begäran i ljuset av den undersökningen , alltså så snabbt som möjligt efter att undersökningen slutförts .
exceptionellt finansiellt stöd till kosovo
nästa punkt på föredragningslistan är betänkande ( a5-0022 / 2000 ) av brok för utskottet för utrikesfrågor , mänskliga rättigheter , gemensam säkerhet och försvarspolitik om rådets förslag till beslut om exceptionellt finansiellt stöd till kosovo ( kom ( 1999 ) 0598 - c5-0045 / 00 - 1999 / 0240 ( cns ) ) .
jag har fått veta att vår föredragande är försenad några minuter .
jag föreslår att vi inleder debatten omedelbart .
föredraganden är på väg hit och kommer att tala så fort han anlänt .
jag lämnar därför ordet till bourlanges i hans egenskap av föredragande av yttrandet från budgetutskottet .
herr talman ! denna fråga är viktig och brådskande och parlamentet , som ombetts av kommissionen att snabbt uttala sig , gör det också , för man skall veta att i dag dör män och kvinnor i kosovo , helt enkelt för att det är 25 grader kallt , att dessa människor utför ett enormt arbete för att garantera ett minimum av underhåll och att de inte får betalt .
vi har därför mottagit en begäran om brådskande förfarande som vi beviljar .
man ber oss om 35 miljoner euro .
vi är överens om att ge ut dem och vi ber kommissionen att visa prov på stor vaksamhet så att beloppen verkligen betalas ut så fort som möjligt när beslutet väl har fattats .
det är fråga om makroekonomiskt stöd .
det orsakar reaktioner på vissa ställen eftersom de liberala idealen inte respekteras som består i att ingripa ekonomiskt för att stödja en administration .
vår uppfattning är att det är grundläggande att bidra till att inrätta en administration i kosovo och att det inte alls är absurt att direkt bidra till att betala de offentliga tjänstemännen i denna region .
det skulle för övrigt ha varit något mycket användbart som vi skulle ha kunnat göra i ryssland under hela 90-talet för att undvika denna stats upplösning .
det andra stora problemet är att man vänt sig till oss , givarna har gjort åtaganden men vi är uppenbarligen de enda som betalar .
de andra betalar inte .
vi kräver att denna unilaterala situation skall upphöra när det gäller att begära ekonomisk hjälp .
vi önskar att kommissionen gör utfästelser när det gäller våra ändringsförslag i det hänseendet .
vi vill knyta beviljandet av hela stödet till mobiliseringen av pengar som övriga givare är skyldiga .
inte för att begränsa , för att knussla med vårt ekonomiska stöd till kosovo utan tvärtom för att se till att vårt stöd kommer utöver det från övriga givare .
ur den synvinkeln är den bestämmelse som föreslås en bestämmelse om stöd i två etapper och den andra bör frigöras när givarna visat att de är intresserade .
avslutningsvis ställer vi tre frågor till kommissionen i detta hänseende : för det första måste den på ett regelbundet sätt ge oss förteckningen och beloppen när det gäller bidrag från övriga givare .
vi vill veta vad de övriga betalar när vi betalar .
för det andra vill vi ha en exakt lägesrapport över anbudsinfordran och deras åtagandetakt .
man sade oss under budgetförfarandet att det var brådskande att rösta för pengarna till kosovo och enligt den information vi förfogar över har hittills ingen anbudsinfordran offentliggjorts eller inletts .
det är allvarligt eftersom det försenar hela återuppbyggnaden av kosovo .
avslutningsvis , och det är konsekvensen av vad jag just sagt , vill vi att kommissionen mycket regelbundet , varje månad , informerar budgetutskottet om läget för verkställandet av utgifterna .
vi har papper från kommissionen där man talar om bestämda åtaganden .
vi behöver inga bestämda åtaganden , vi behöver åtaganden helt enkelt och vi behöver veta vad som verkligen betalats och framför allt vad som inte betalats .
kosovo har lidit alltför mycket av försenade betalningar .
herr talman ! när vi i dag talar om kosovo , vilket vi ju ofta har gjort , bör vi också någon gång avlägga räkenskap om vad som redan har gjorts i kosovo , eller om det över huvud taget redan gjorts något .
jag anser att man redan har tagit några små steg på vägen mot en normalitet , och man skulle åtminstone vilja räkna upp dem inom ramen för en sådan debatt .
det finns från och med den 9 februari ett s.k. interimsråd - man kallar det kosovo transitional council - , där både de politiska partierna , minoriteterna och the civil society är representerade , och som skall fungera ungefär som ett interimsparlament .
det är bra , det välkomnar vi , men jag tror att man också måste ge dem ett instrument i handen och en strategiplanering för det som de egentligen bör förbereda , ty i höst planerar man att hålla val .
ingen vet riktigt vad dessa val skall leda till , och vilket parlament som skall bildas .
ingen vet vilka befogenheter detta parlament sedan skall ha gentemot unmik .
det betyder att det finns många svårbedömbara saker som vi inte informeras om och som andra förmodligen inte heller kan riktigt förstå .
just albanerna , som nu integreras i detta interimsråd , borde egentligen få en något bättre uppfattning om vad som väntar dem .
vid sidan av det ekonomiska arbetet , vid sidan av återuppbyggnaden , måste man ovillkorligen också tänka på hur man skall åstadkomma någon samexistens mellan serber , albaner och andra minoriteter - exempelvis också zigenarna - så att det , på vägen till samexistens , någon gång i en nära framtid förhoppningsvis kan äga rum en försoning .
jag vill än en gång räkna upp vad det redan finns av faktiska saker som vi kan glädja oss åt .
när det gäller förvaltningen finns det nu 34 skatteinspektörer .
människorna uppmanas nu också att betala sina skatter även där , ty på sikt kan det ju inte gå an att alla bara är beroende av eu : s och andra givares portmonnäer ; en del måste man även på detta område åstadkomma på egen hand .
det kan dessutom fastslås att av 19 departement har redan 4 en administrativ ledning , vilket också är ett framsteg jämfört med vad vi tidigare haft där .
vi har dessutom något som är mycket viktigt för den rättsstat som vi ju vill bygga upp .
vi har 130 domare och åklagare , som nu har avlagt eden , och som kan ta upp sitt arbete för att skipa rätt , för att också litet grand berika toleranskulturen där en aning och naturligtvis också åtminstone komma förbrytelserna på spåren och då också kunna döma .
det som också är bra , det vill jag erinra om , är det faktum att den gamla uck nu är integrerad i återuppbyggnaden av detta land .
jag ansluter mig helt och fullt till det som budgetutskottet har sagt i fråga om finansieringen , och jag anser att vi måste erinra kommissionen om att den verkligen måste insistera på att andra givare äntligen betalar sin andel .
eu-kommissionen kan inte betala för allting .
den är där nere ansvarig för återuppbyggnaden , den är ansvarig för den fjärde pelaren , men den kan inte också alltid betala kouchners löpande kostnader .
det kan man göra en eller ett par gånger , men jag tror att fn : s givare också måste bidra till det , och där finns det ett mycket stort hål , som inte är fyllt , och som vi inte kan fylla .
vi har en stor uppgift i återuppbyggnaden , det är vår uppgift , och vi bedöms efter hur vi utför denna uppgift !
herr talman ! jag vill göra några preciseringar .
risken i en debatt är alltid att vi som medverkar upprepar oss för mycket .
men jag skall koncentrera mig på fyra punkter .
till att börja med vill jag fastslå att unionen är den största bidragsgivaren till återuppbyggnaden av kosovo .
och till albright kan jag säga att detta har stått i tidningen på senare tid , och siffrorna ljuger inte .
detta råder det ingen tvekan om , även om man kunde önska att det inte vore fallet .
unionen har beslutat att bidra med ytterligare 35 miljoner euro i makrofinansiellt stöd till återuppbyggandet av kosovo , mot bakgrund av en rapport från fmi där man uppskattar att återuppbyggandet kräver ytterligare 115 miljoner .
jag vill nämna för pack att jag med henne är helt överens om att kommissionen måste uppmana de övriga bidragsgivarna att uppfylla sina löften .
dessutom vill jag ge uttryck för min oro - en mycket stark sådan - över vissa ministrars uttalanden på det senaste ekofin-rådet , som visar att man vill att en av det portugisiska ordförandeskapets prioriteringar skall vara att den budgetplan som man enades om i berlin under inga omständigheter ändras .
detta innebär ett ifrågasättande av det avtal som parlamentet med stora svårigheter lyckades uppnå med rådet i december , enligt vilket man , när kommissionen lägger fram ett flerårigt program för återuppbyggandet , skall vidta en granskning av budgetplanen .
därför vill jag uppmana dessa ministrar att inte ifrågasätta det avtal som var så svårt att uppnå .
jag vill be kommissionen , och det gläder mig att kommissionär solbes är här i kväll , att i god tid lägga fram detta fleråriga finansieringsprogram , med tillhörande rapport , enligt parlamentets begäran , så att det kan beaktas i framtagandet av budgetförslaget till nästa budget , i överensstämmelse med det som vi har blivit lovade .
slutligen vill jag poängtera att vi även om vi nu har kommit överens om 35 miljoner , vet att det bara är en droppe i havet och att det inte är tillräckligt , och därför måste vi så snart som möjligt uppnå en överenskommelse om ett flerårigt program för det så nödvändiga återuppbyggandet av kosovo .
herr talman , kolleger ! jag ber er ursäkta att jag är försenad , men i dag är tyvärr denna andra politiska fråga fortfarande på föredragningslistan .
utskottet för utrikesfrågor , mänskliga rättigheter , gemensam säkerhet och försvarspolitik rekommenderar att ni lösgör dessa 35 miljoner euro , och den rekommendationen ger man eftersom dessa pengar verkligen kan komma de drabbade människorna till godo .
det vi är kritiska till är inte så graverande att vi inte vill hjälpa människorna där nere .
men det betyder inte att vi glömmer bort kritiken .
vi skulle naturligtvis redan ha kommit mycket längre i vårt förfarande om rådets förvaltning inte hade glömt bort att på ett tidigt stadium informera europaparlamentet och officiellt lämna information till det .
endast på så sätt hade vi kunnat genomföra ett verkligt förnuftigt , djupgående samråd i saken .
jag ber förvaltningen att se till att detta inte kan hända i framtiden .
endast för de drabbade människornas skull är vi beredda att bortse från det och dra konsekvenserna av det .
men vi måste se till att vi här inför bestämda villkor .
ett villkor är att pengarna ges dit där de kommer att användas på ett klokt sätt , och inte till dem som möjligen kan använda pengarna för att tjäna andra syften , dvs. dessa pengar bör verkligen gå in i kouchners ansvarsområde och inte till andra områden .
för det andra : även om kommissionen och rådet här intar en annan ståndpunkt , eftersom de där ser realistiska problem , anser vi att de andra givarna också måste uppfylla de åtaganden som de har ingått .
detta är en mission som står under fn : s ansvarsområde , och det får inte vara så att enbart europeiska unionen uppfyller sina förpliktelser !
de andra givarländerna måste uppfylla sina förpliktelser på samma sätt under denna tidsrymd till gagn för de drabbade människorna .
detta får mig att anse att vi i framtiden rent allmänt måste befatta oss mycket intensivare med denna fråga , och inte bara när det gäller detta konkreta projekt , utan hela utvecklingen i sydosteuropa , och den hjälp som lämnas där .
detta är återigen ett exempel för att europeiska unionen är beredd att hjälpa till att ge pengar , men att den politiska ledningen inte är enhetlig .
vi har så många samordnare , som är ansvariga inför så många arbetsgivare , att vi snart måste tillsätta en samordnare för samordnarna .
men det kanske vore bättre om de ansvariga instanserna i europeiska unionen och de andra institutionerna , från osse till förenta nationerna - skulle sätta sig ned för att införa ett enhetligt , samordnat förfarande , och granska hur man verkligen kan hjälpa människorna där .
jag vet att man inom kommissionen intensivt funderar över hur man skall uppnå detta , men om europeiska unionen bidrar med den största delen , då skall den också ha hand om ledningen där och sedan sköta det på ett enhetligt sätt , så att människorna verkligen blir hjälpta .
det är ingen mening med att vi här snarast har en konkurrens mellan de olika internationella inrättningarna och sammanslutningarna , i stället för att kraften verkligen utnyttjas för att hjälpa människorna på platsen !
när jag ser att givarkonferensen för stabilitetspakten hela tiden skjuts upp , nu till slutet av mars , och att ingen vet vilka projekt som verkligen ligger bakom , när man inte kan överblicka på vilket vis det verkligen kan genomföras , och det hela tiden ges nya presskonferenser , då verkar detta inte vara rätt sätt att skapa fred och försoning mellan människorna i denna del av europa !
av den anledningen , kära kommission , kära ordförandeskap i rådet , vill vi också ta detta till anledning för att uppmana er att gripa detta politiska initiativ , så att vi inte åter hamnar i en sådan nödsituation att vi i slutet av en månad måste ordna upp betalningsförmågan , utan att det därmed kan ställas upp en långfristig strategi för hjälpen i denna region , och jag hoppas att ni då äntligen kan uppfylla era politiska förpliktelser , och att det inte fortsätter så som vi har upplevt det under de senaste månaderna !
herr talman ! när alliansen engagerade sig i kosovo var det med målsättningen att i denna provins återupprätta villkor som gör det möjligt för dem som så vill att stanna kvar , återvända till sina rötter och till sin egen kultur .
om alliansen i dag är närvarande på fältet är det med samma målsättning .
i förrgår lyssnade jag med tillfredsställelse till en intervju med en befälhavare i kfor som berättade att saker och ting började fungera bättre i kosovo och att normerna för brottsligheten återgått till en acceptabel nivå , framför allt när det gäller säkerhet .
de som befinner sig på fältet för att företräda europa och fortsätta med dessa målsättningar , och jag tänker särskilt på den särskilda representanten för förenta nationernas generalsekreterare , är nära att ge upp , just på grund av det faktum att situationen förbättrats och man talar mindre om kosovo , och att det därför är mindre uppenbart hur brådskande hjälpen är som behöver beviljas .
vi måste arbeta för att se till att epoken med kommers ersätter den med krigsherrarna , i denna provins liksom i hela balkan i allmänhet .
det ekonomiska stödet är i det hänseendet en beståndsdel som förvisso är grundläggande när det gäller möjligheter till åtgärder för dem som befinner sig på fältet .
jag upprepar här doris packs uttalande och jag betonar att vi i europaparlamentet måste ta vårt ansvar i detta hänseende , men vi skall naturligtvis se till att vi inte är ensamma om det .
herr talman , herr kommissionär , mina damer och herrar ! först vill jag tacka föredraganden , kollegan brok , så hjärtligt för hans betänkande .
om rådet hade arbetat så snabbt som kollegan brok gjort , då skulle vi i själva verket ha kommit mycket längre .
rådets försummelse kan man här verkligen beklaga !
föredraganden och betänkandet utgår helt riktigt från att vi bör och måste lämna snabb hjälp , men de utgår också helt riktigt från att vi inte skall lämna obegränsad eller godtycklig hjälp .
här vill jag i synnerhet hänvisa till ändringsförslag 5 , där det helt klart fastslås att man med hjälp av medlen från det särskilda ekonomiska stödet uteslutande kan och får finansiera sådana budgetbehov i kosovo , som uppstår i offentliga / halvoffentliga , kommunala och övriga förvaltningar och institutioner , som direkt eller indirekt kontrolleras av unmik .
det måste stå klart , herr kommissionär , att vi stöder unmik , vi stöder de institutioner som inrättats av förenta nationerna , i synnerhet naturligtvis pelare 4 , och det går inte an att vi stöder parallella strukturer som har bildats i kosovo och fortfarande finns kvar där .
vad skall nu göras med dessa pengar ?
jag vill särskilt hänvisa till de mänskliga rättigheterna .
västmakterna har i kosovo kämpat för de mänskliga rättigheterna .
vad sker i dag i kosovo ? den stora aktionen för att driva bort serberna kunde stoppas , men nästan dagligen sker det oacceptabla saker , människor dödas , människor hindras att leva där , och att leva på sitt vis .
dagligen sker det angrepp på serber , på zigenare , på bosnier , men det sker också fortfarande angrepp på albaner .
jag blev förskräckt när jag läste betänkandet , om det nu stämmer att en albansk läkare , som säkerligen med stora svårigheter arbetat i sjukhuset i mitrovic i den serbiska delen , slutligen gav upp att arbeta för sin befolkning i detta sjukhus , eftersom han hela tiden hotades till livet .
detta är händelser och situationer som vi inte kan acceptera .
jag har hört - om det stämmer vet jag inte - att serberna fortfarande rent av driver en gruva i kosovo , i den serbiska delen .
det finns åtminstone rykten om att serbisk milis fortfarande är aktiv .
för mig är det betydelselöst om det är en serb , en zigenare , en bosnier eller en alban som hotas eller dödas i kosovo .
för mig är det betydelselöst vem som arbetar på att dela kosovo .
det som är avgörande för mig är att de organ som finansieras av oss uppnår det som vi vill uppnå , nämligen ett multietniskt kosovo , ett liv sida vid sida i kosovo .
vi behöver mer polis , det finns absolut inte tillräckligt med polis .
vi behöver ett oberoende rättsväsende - det är säkert svårt att bygga upp - och vi behöver också anslag för den höge kommissionären för de mänskliga rättigheterna .
allt detta måste ske , och det måste ske snabbt .
om vi inte snabbt lämnar hjälp , då kommer situationen att förvärras , och det kan uppstå nya konflikter och krissituationer .
därför anser jag att det var rätt att vi handlade snabbt , att vi bekräftade att det var brådskande , och att vi ställer pengarna till förfogande .
men vi vill se vad som görs , och vi vill också se resultat i kosovo , och jag ber kommissionen att se till att dessa pengar också används med framgång , i synnerhet för att bygga ut polisväsendet och rättsväsendet .
- herr talman !
till en början ett stort tack till ledamöterna , och i synnerhet till föredraganden , för den snabba behandlingen av denna fråga .
det kommer utan tvivel göra det möjligt för oss att snabbt frigöra medel till kosovo och ta oss an de orosmoment som både swoboda och pack har påtalat .
i den här kvällens debatt tycker jag mig märka tre starka orosmoment .
för det första är det sant att vi , även om det har skett stora framsteg , och där kan nämnas tullförvaltningen , bankförvaltningen och skatteförvaltningen , måste fortsätta framåt .
framåt mot en finansiering av vad ?
där har vi den första punkten där det råder en viss oenighet .
ni föreslår i ett av era ändringsförslag att enheterna som är föremål för unionens finansieringsbidrag skall begränsas mer . till exempel i ändringsförslag 3 och 5 .
emellertid bör man , enligt vår uppfattning , i båda avseendena lämna större handlingsutrymme åt förenta nationernas förvaltning som känner till förhållandena på platsen bättre än vi .
vi anser att det skulle innebära stora praktiska svårigheter att redan på förhand definiera vart resurserna skall gå .
vi måste utan att tveka förlita oss på dem som där på plats , på ett bättre sätt än vi , kan fatta vissa beslut .
det andra orosmoment som jag har förstått att vissa av er känner av - det lades till att börja med fram av bourlanges , och det har upprepats av andra - gäller det som händer med övriga bidragsgivare .
är det så att kommissionen gör en överdriven insats , medan de övriga struntar i att samarbeta ?
vissa av ändringsförslagen i ert betänkande pekar i den riktningen .
till exempel ändringsförslag 1,2 och 4 .
jag kan tala om för bourlanges och för dem som har lagt fram denna fråga , att det främsta problemet inte gäller tanken som sådan , som vi är helt eniga i .
det främsta problemet är att fördelningen av bördan mellan de olika bidragsgivarna för närvarande har fastställts - och det är sant - i uttalandena av high level steering group , men det stämmer också att de saknar juridiskt värde , att det endast rör sig om ett politiskt åtagande .
det är anledningen till att vi ber att ändringsförslag 1 , och vi har meddelat brok detta , med bibehållen andemening skall formuleras på ett annat sätt så att det inte innehåller några villkor för tilldelningen av gemenskapens resurser .
det samma gäller ändringsförslag 2 , som vi också finner godtagbart om det bara justeras något , eftersom vi anser att idén vad det finansiella stödet beträffar i sig är korrekt .
ungefär samma sak gäller ändringsförslag 4 .
i denna konkreta fråga är det möjligt att vi har ett mer positivt besked till bourlanges .
rådet är redan vidtalat , så att det skall låta sitt beslut omfatta ett uttalande av kommissionen där detta villkor fastslås .
det vi föreslår är närmare bestämt , vad det andra bidraget beträffar , att det exakta totalbeloppet och tidpunkten för den andra delutbetalningen skall avgöras med hänsyn till kosovos externa finansiella behov och stödet från övriga bilaterala bidragsgivare .
vi fastslår med andra ord inget villkor , eller vi tror att det är mer effektivt att inte fastslå något villkor från början , och ändå gör vi det beträffande detta eventuella frigörande av den andra delutbetalningen .
på det viset kommer vi inte att ha några problem med att agera omedelbart , vi skapar inga problem för befolkningen i kosovo , men däremot tvingar vi de övriga bidragsgivarna att genomföra sina finansiella insatser på samma sätt som vi gör .
ett tredje problem har påtalats av dührkop beträffande de fleråriga programmen .
jag kan påminna om att projekten är fleråriga .
i programmen måste man givetvis ta hänsyn till det årliga budgetstödet .
till slut vill jag kommentera de önskemål som har framförts om ytterligare information .
å ena sidan har man bett oss underlätta utvecklingen av anbudsförfarandet för parlamentet , och på den punkten kan jag tala om för er att kommissionen redan förra veckan hade tillfälle att ge parlamentets budgetutskott en lägesrapport om de kontrakt och betalningar som har utförts sedan task force började fungera i kosovo .
kommissionen kan lova att även framöver regelbundet informera parlamentet om de anbudsförfaranden som offentliggörs .
vår önskan är att detta även läggs ut på internet , så att största möjliga insyn ges i denna konkreta fråga .
en annan sak jag vill kommentera är övrig information som kan vara av betydelse för parlamentet vad gäller det makroekonomiska stödet .
i det avseendet kan jag även meddela att kommissionen är villig att regelbundet informera ordförandena i de olika parlamentsutskott som är involverade i frågan , under konfidentiella former om den information som ges förutsätter detta , samt utifrån de olika planer som tillämpas för de makroekonomiska stödåtgärderna .
ett stort tack till alla ledamöter , och jag hoppas att vi i och med rådets slutgiltiga beslut kan få loss dessa medel och förverkliga ett positivt stöd som gör det möjligt för oss att fortsätta med de viktiga insatser som görs i kosovo från olika håll för att uppnå den situation som vi alla önskar med en ökad förståelse och fred .
herr talman ! jag gläds åt att åsikterna från parlamentet , särskilt budgetutskottet , och kommissionen är så samstämmiga , och vi försäkrar att för vår del kommer vi alltid att troget hjälpa kommissionen att genomföra sin uppgift .
jag känner ändå en viss oro när jag lyssnar till kommissionären jämfört med de åtaganden som gjorts av enheterna inom budgetutskottet .
det beslutades tydligt - jag säger inte att det var bra eller dåligt , men det var ett avtal - det beslutades tydligt mellan kommissionens enheter och budgetutskottet att man var överens om ändringsförslag 4 och 7 , dvs. man var överens om idén att knyta mobiliseringen , genomförandet , av den andra delen av det makroekonomiska stödet till respekten för de åtaganden som tidigare gjorts av givarna .
men jag tyckte mig förstå när jag lyssnade till solbes att detta åtagande skulle ske på ett diskret sätt .
herr kommissionär ! ett avtal är ett avtal .
ja eller nej , bekräftar ni det godkännande som gjorts av era enheter i budgetutskottet eller släpper ni detta villkorande , vilket skulle innebära att ni bryter ett åtagande mot oss ?
. ( fr ) nej , herr bourlanges , jag tror att det handlar om ett sakproblem .
problemet är : hur skall vi styra den kompromiss vi accepterat .
vad jag föreslog er , vad jag säger igen , är att kommissionen skall göra ett uttalande , i rådets beslut , i följande riktning :
det exakta beloppet och tidpunkten för att inleda den andra delen kommer i sinom tid att beslutas med hänsyn till utvecklingen av kosovos yttre ekonomiska behov och bidrag från andra bilaterala givare .
därför anser vi att vi fullständigt respekterar det som vi kommit överens om .
jag begär bara att kommissionen skall informera budgetutskottet innan den andra delen genomförs .
( fr ) jag instämmer helt , och det kommer vi att göra .
altener
nästa punkt på föredragningslistan är betänkande ( a5-0011 / 2000 ) av langen om förlikningskommitténs gemensamma utkast till parlamentets och rådets beslut om ett flerårigt program för främjande av förnybara energikällor inom gemenskapen - altener ( c5-0333 / 1999 - 1997 / 0370 ( cod ) )
herr talman ! jag tackar langen - även om han inte själv är närvarande här - för det arbete som han lagt ner för att driva igenom programmet såväl i parlamentet som i rådet .
projektet har varit långvarigt och besvärligt .
man måste även i fortsättningen satsa särskilt mycket på sådan forskning som kartlägger användningen av förnybara energikällor .
även om det nya direktivet innehåller mycket gott är det dock också behäftat med brister .
ett exempel på detta är torven .
torv får inte placeras i samma grupp som fossila bränslen .
kan man inte direkt klassificera torven som en förnybar , icke-fossil energikälla måste man särskilt med tanke på miljöbeskattningen definiera en egen klass för den .
det är inte rättvist att torven värderas på samma sätt som exempelvis stenkolen .
utvecklingen av förnybara energikällor är en dellösning för att avskaffa unionens beroende av importerad energi .
forskningen är av speciellt stor betydelse också med tanke på eu : s nästa utvidgningsrunda .
beroendet av importerad energi berör allra värst just flera östeuropeiska länder vars ekonomiska struktur fortfarande lider av det beroende av rysk energi som skapades under sovjettiden .
eu måste hålla fast vid kyotos klimatprotokoll .
vi är ju alla bekymrade över miljön och våra barns framtid .
de förnybara energikällornas andel av den totala energiproduktionen måste ökas , men det måste också göras med förnuft .
vi måste komma ihåg att vi inte på länge än kan bygga vår grundläggande energiproduktion på förnybara energikällor .
där behövs energi som skonar klimatet , kärnkraft .
herr talman ! å pse-gruppens vägnar är jag positiv till att vi har kommit fram till ett resultat i förlikningsförfarandet beträffande altener ii-programmet .
men först vill jag tacka föredraganden , kollegan langen , för hans verkligt bra arbete med detta betänkande .
jag vill också tacka ledaren för delegationen till förlikningskommittén , kollegan provan .
ty som langen just sade var det verkligen en hård kamp i förlikningskommittén .
men vi kan i dag se att resultatet av förlikningen också absolut mycket tydligt visar vad europaparlamentet förmår .
langen påpekade att en rad punkter beträffande innehållet och krav från parlamentet införlivats , och när det gällde den viktigaste konflikten med rådet , anslagen till detta fleråriga program för att främja de förnybara energikällorna i gemenskapen , kunde vi - det har redan sagts - enas med rådet någonstans på mitten .
det är inte tillfredsställande , det vill jag också säga helt klart .
men vi har gått med på denna kompromiss , eftersom det var viktigt för oss att detta program nu verkligen kan startas mycket snabbt .
ty under de närmaste åren skall andelen förnybara energikällor fördubblas till minst 12 procents andel av energiförbrukningen .
det är europeiska unionens uttalade mål .
där har altener-programmet verkligen en nyckelroll , som enda eu-program med den uteslutande målsättningen att främja förnybara energikällor .
med detta nya femårsprogram måste dels åtgärderna från altener i-programmet utökas .
hit hör bland annat fördjupningen av informations- och erfarenhetsutbytet mellan aktörerna på området med alternativa energikällor , bland annat utbyggnad av lokala och regionala energiagenturer , uppbyggnad av nya nät och stöd till bestående nät . detta är bara några exempel .
men det som är särskilt viktigt när det gäller altener ii-programmet är - anser jag - de nya åtgärderna för att underlätta att de förnybara energikällorna får genomslagskraft på marknaden , och de nya åtgärderna för att genomföra , åtfölja och övervaka gemenskapens strategi och gemenskapens åtgärdsplan .
det föreligger nu ett arbetsdokument från kommissionens enhet rörande en kampanj för ett genombrott , vilken ju är en väsentlig beståndsdel i denna gemenskapsstrategi .
det som här planeras är stöd på alla väsentliga områden i fråga om förnybara energikällor .
detta altener-program måste verkligen åtfölja och stödja denna kampanj .
de totala investeringskostnaderna för kampanjen har beräknats till ca 30 miljarder euro .
därav skall 75 - 80 procent komma från privata källor , och härtill kommer allmänna medel från medlemsstater och regioner .
här kan altener-programmet ge viktiga nya impulser för investeringar , underlätta dem och hjälpa oss så att vi verkligen kan uppnå vårt mål beträffande miljöskydd , ekonomi och nya arbetstillfällen .
herr talman , fru kommissionär ! även jag vill tacka langen för det goda arbete han lagt ned i detta viktiga ämne .
det slutresultat av förlikningen avseende altener-programmet som förlikningskommittén lagt fram är efter ett antal svåra turer åtminstone nöjaktigt .
största delen av parlamentets ändringsförslag har beaktats , och som en positiv sak måste man konstatera att finansieringsbeloppet för programmet höjts till 77 miljoner euro .
när det gäller ökad användning av förnybara energikällor har unionen ambitiösa mål .
i förhållande till dessa mål är anslaget emellertid mycket litet .
det måste användas till pilotprojekt , forskning , informationsutbyte samt till att bilda positiv opinion för användningen av förnybara energikällor .
huvudansvaret för att öka användningen av förnybara energikällor vilar på medlemsstaternas axlar .
förhoppningsvis väcker detta program medlemsstaterna till att bedriva en beslutsam verksamhet för att öka användningen av förnybara energikällor .
men även unionen måste i framtiden öka sin egen satsning för att främja användningen av förnybara energikällor och se till att den förnybara energin utan hinder kan komma in på marknaden .
att främja användningen av förnybara energikällor är särskilt viktigt med tanke på miljön .
de förnybara energikällorna minskar beroendet av importerad energi och ökad användning av dem förbättrar konkurrenskraften .
europa kan också uppnå en ledande position inom den industri som levererar de utrustningar som behövs för att använda förnybar energi .
man måste också komma ihåg att användningen av förnybara energikällor har en positiv inverkan på den regionala utvecklingen och sysselsättningen .
även jag vågar nämna torven .
torven finns inte med på listan över förnybara energikällor .
den är dock åtminstone i finland en viktig , långsamt förnybar energikälla som används på ett hållbart sätt .
jag hoppas att den i framtiden kan tas med på listan över förnybara energikällor .
fru kommissionär , kära kolleger ! gruppen de gröna gläds åt den överenskommelse som gjorts och vårt tack går till alla dem som förhandlat så bra för ett ändringsförslag som de gröna nästan var upphovsmän till .
det är intressant för mig , som är ny här i parlamentet , att konstatera att man i budgeten planerar för hundratals miljoner euro per år för tobaksodling .
det är en begränsad sektor av ekonomin som nästan inte skapar någon sysselsättning , som inte är konkurrenskraftig på världsnivå .
jämfört med detta konstaterar jag de summor som står på spel för förnybar energi som inte bara är en ekologisk beståndsdel utan också är förutbestämd att få en avsevärd ekonomisk uppgång .
när man ser de marknadsandelar som små länder såsom danmark lyckats förvärva på detta område , tack vare att de var de första på marknaden , tror jag det manar till eftertanke och att vi på lång sikt verkligen måste öka budgeten för förnybar energi .
ett sista ord när det gäller programmet : jag tror att det är mycket viktigt att de förnybara energikällorna , om de skall kunna utvecklas på lång sikt , är förankrade i regionerna där de kan bidra till ekonomin och till att skapa sysselsättning .
om 50 procent eller mer av energimixen skall kunna komma från förnybara energikällor kan man inte nöja sig med vissa hot spots som på kort sikt blir mer lönsamma .
herr talman ! jag vill inleda med att gratulera herr langen för hans arbete .
aktiviteterna inom ramen för altener-programmet kommer att främja förnybara energikällor och jag anser att sådana program förtjänar finansieringsstöd på utvecklingsstadiet då de erbjuder enorma kommersiella möjligheter i framtiden .
av detta skäl är jag särskilt glad att se att pengarna satsats på små och medelstora företags projekt .
de internationellt överenskomna målen för minskade utsläpp kan inte uppnås genom dessa program enbart .
i detta hänseende måste man komma ihåg att energipolitiken förblir inom ramen för nationella befogenheter .
det är ytterst viktigt att de nationella regeringarna ger sitt fulla stöd för att få en effektivare energianvändning och för att utveckla förnybara energikällor .
jag är förtjust över att irland nyligen meddelade att man där kommer att använda 125 miljoner irländska pund för att utveckla en miljömässigt hållbar energisektor .
jag hoppas att altener-programmet skall medverka och leda till fler initiativ .
såsom korrekt fastslås i den slutgiltiga texten kan åtgärder som dessa spela en roll för att minska regionala skillnader .
jag kan intyga att jag redan har mottagit bevis på stort intresse för altener-programmet från min egen valkrets leinster , en region som till en betydande del ligger inom irlands enda mål 1-region .
jag stöder alla insatser för att minska klyftan inom ekonomisk utveckling av infrastrukturbestämmelser , inklusive energisektorn .
kort sagt , vi står inför en stor utmaning för att klara av våra åtaganden att begränsa utsläppen av växthusgaser från energisektorn enligt kyoto-protokollet medan vi samtidigt främjar tillväxten i våra ekonomier .
altener-programmet skall vara ett värdefullt bidrag till medlemsstaternas samlade insatser .
- herr talman , mina damer och herrar !
jag vill börja med att uttrycka min glädje över den överenskommelse som har uppnåtts angående programmet altener ii i förlikningskommittén och ansluta mig till de uttalanden som har gjorts av tidigare talare , och givetvis påpeka att denna överenskommelse kommer att innebära att programmet altener inom kort tas med i ramprogrammet för energi .
allt detta kommer att leda till en ökad samordning , insyn och effektivitet i våra energiprogram , i vilka även programmet save måste införlivas , vilket vi snart kommer att diskutera .
jag anser att parlamentets arbeten under den här perioden har hållit hög standard , och därför gratulerar jag föredragande langen och även de olika talare som har hållit anföranden , både i kommissionen och här i parlamentet .
det är uppenbart att det har förts diskussioner , vi blev tvungna att söka förlikning , precis som föredraganden och caudron påpekade för en stund sedan , för under det första mötet uppnåddes inga resultat , och man blev därför tvungen att samlas en andra gång , trots att siffrorna inte heller var överdrivet höga .
men jag anser att vi till slut lyckades uppnå ett rimligt avtal som i likhet med alla avtal inte är fulländat , men som jag tror gör det möjligt att fortsätta med de projekt som vi hade på gång .
därför vill jag upprepa mina gratulationer till föredraganden langen för det arbete han har utfört , tacka alla talare och naturligtvis lovorda vice ordförande provans agerande under förlikningsförfarandet som i stor mån bidrog till att uppnå ett positivt resultat .
jag vill även lovorda rådets förnuftiga och flexibla attityd .
save
nästa punkt på föredragningslistan är betänkande ( a5-0010 / 2000 ) av ahern för europaparlamentets delegation till förlikningskommittén om förlikningskommitténs gemensamma utkast till europaparlamentets och rådets beslut om att anta ett flerårigt program för att främja en effektiv energianvändning - save ( c5-0334 / 1999 - 1997 / 0371 ( cod ) ) .
. - ( en ) fru talman ! jag vill tacka rådet och kommissionen för ett bra och omsorgsfullt förlikningsförfarande där alla var vid gott humör vilket inte alltid är fallet .
det är ett nöje för mig att säga att jag anser slutresultatet av förlikningen som mycket tillfredsställande för parlamentet då den gemensamma texten innehöll alla dess ändringsförslag antingen hela texten eller i omformulerad form .
det belopp som slutligen anslogs till programmet är också en betydande förbättring mot rådets förslag vid den andra behandlingen som vi ansåg som helt oacceptabelt och vi har lyckats få betydande framgång där .
jag föreslår därför att denna kammare antar förslagen för save-programmet och slutsatsen vid förlikningen vid tredje behandlingen .
jag vill påminna kammaren om att vid andra behandlingen godkände parlamentet detta betänkande innehållande åtta ändringsförslag , inklusive ett återinförande av kommissionens ursprungliga budget .
kommissionen godkände fem av de föreslagna ändringsförslagen , inklusive budgetanslaget , och jag tackar kommissionen för deras fortsatta stöd om budgeten under förlikningsförfarandet då det som rådet hade föreslagit var oacceptabelt .
under förfarandet kom man överens om vilka undersökningar och insatser som skulle planeras , genomföras , kompletteras och utvärdera gemenskapsinsatserna .
kompromissformuleringar enades man om för fem andra ändringsförslag inklusive lagstiftnings- och icke lagstiftningsåtgärder och inrättandet av lokala energicentra och , något mycket viktigt , energikontrollsystem en som skall följa upp utvecklingen av ökad energieffektivitet .
jag hoppas att ni alla skall hålla med om att detta är en viktig utveckling .
frågan om det finansiella anslaget försvarades hårdnackat av parlamentet ställt mot rådets mycket låga öppningserbjudande .
i varje fall fick vi lova att hålla flera sammanträden innan rådet slutligen höjde beloppet avsevärt .
vi fick en ökning med 2 miljoner mot deras första förslag , vilket var en betydande höjning som jag kan rekommendera er och som kommissionen bekräftade skulle räcka för att den skulle kunna genomföra programmen .
detta var ett viktigt ställningstagande för oss .
jag skulle dock vilja framföra att det är och har alltid varit en mycket blygsam budget och därför är finansieringen för detta program mer symbolisk än reell .
finansieringen för att spara energi görs fortfarande huvudsakligen av medlemsstaterna .
vi måste komma ihåg det när vi godkänner detta program .
om det är fråga om mer symbolism än realitet i fråga om det som vi kan uppnå på gemenskapsnivå är det synd för det finns mycket entusiasm på lokal nivå för åtgärder , däribland gemenskapsåtgärder , för energibesparing .
ett område där gemenskapen kan hjälpa till är att skapa kontakter mellan lokala aktörer så att de inte behöver starta om från början i varje region .
vi har en betydelsefull roll att spela i gemenskapen inom europeiska unionen i detta avseende .
save är det enda program som täcker hela gemenskapen och som är avsett att främja en rationell energianvändning .
det är inriktat på icke tekniska områden för att skapa energieffektiva infrastrukturer och ändamålet med programmet är att skapa en miljö för att främja investeringar och en effektiv energianvändning .
här behöver vi inse att det även finns en marknadsmöjlighet inom industrin för energibesparingar .
vi har hört en massa om konkurrenssvårigheter inom förnybara energikällor men energieffektivitet sparar pengar för företag , sparar pengar överallt i själva verket , och därför bör det inte finnas problem här .
det är något som vi alla kan stödja .
jag måste säga , liksom moderskap , även om vi alla stöder det , gör vi ibland mycket lite i det stora hela och rent konkret för att hjälpa mödrar eller människor som är intresserade av energibesparing .
vi kan göra ganska mycket mer med hänsyn till att vi har gjort stora åtaganden för att minska utsläppen av koldioxid och växthusgaser och för att minska beroendet av energiimport .
vi vidtar inte de åtgärder som medborgarna önskar .
vi visar inte på sambandet så att medborgarna verkligen kan göra något konkret i hemmet eller på sina kontor eller i industrin för att stödja åtgärderna mot globala klimatförändringar .
om vi kan föra fram detta budskap skulle det vara en mycket intressant sak att göra .
jag vill återigen tacka alla som hjälpte till i detta förlikningsförfarande .
- fru talman , mina damer och herrar ! jag vill åter igen tacka fru ahern för hennes arbete som föredragande av detta förslag , för hon har i samarbete med övriga parlamentariker bidragit till att man slutligen uppnått ett högst rimligt resultat , som i vissa avseenden även förbättrar en del av kommissionens förslag och naturligtvis det som rådet till en början hade godkänt ur budgetsynpunkt .
precis som ahern så riktigt sade är både budgeten för save- programmet och den för altener-programmet , i första hand symboliska budgetar , för den tyngsta bördan bär länderna , unionens stater , regionerna och även i vissa fall kommunerna .
hur som helst innebär inte dess begränsade volym att den upphör att ha det viktiga symboliska värde som förutsätts av det faktum att det inom gemenskapen som helhet finns en vilja att stödja denna typ av åtgärder som bidrar till att vi verkligen uppfyller våra löften från kyoto och dessutom till att vi uppnår ett större mångfald i våra energikällor , en ökad säkerhet i vår energiförsörjning och , som i fallet med save , att vi närmar oss en lägre konsumtion , ett mer effektivt utnyttjande av energin , och därigenom bidrar till att nå de uppsatta målen .
dessutom står vi nu i samband med dessa program , det vill säga save-programmet för en effektiv energianvändning och altener-programmet för förnybara energikällor , inför en mycket viktig teknisk utmaning , som ur ekonomisk synvinkel kan komma att innebära stora möjligheter för industrin och även för skapandet av sysselsättning i våra länder , och därigenom i hela unionen .
vad beträffar den parlamentariska behandlingen , vill jag upprepa mitt tack till alla de som har agerat och talat , och huvudsakligen föredraganden , för i det förslag som har godkänts av rådet har de flesta av parlamentets ändringsförslag tagits med , praktiskt taget samtliga i det här fallet , om än med vissa ändringar , och jag vill tacka för att man dessutom har lyckats förbättra det första erbjudandet vad medlen beträffar .
det har man lyckats göra med hjälp av nya pengar , så som vi den gången sade , och man har lyckats göra det och samtidigt bevara parlamentets förmåner och behörighet .
från kommissionens sida sett , i detta spel institutionerna emellan , anser jag att det är viktigt , och jag har nöjet att få poängtera detta .
jag vill upprepa mitt tack till alla som har talat , i synnerhet till vice ordförande provan , för hans föredömliga agerande under denna debatt , framför allt under förlikningsprocessen , till ordföranden i utskottet för industrifrågor , utrikeshandel , forskning och energi , och även till föredragande ahern , samt till alla de ledamöter som har deltagit i arbetet .
nästa punkt på föredragningslistan är betänkande ( a5-0009 / 2000 ) av graça moura för europaparlamentets delegation till förlikningskommittén om förlikningskommitténs gemensamma utkast till europaparlamentets och rådets beslut om att inrätta ett enhetligt instrument för finansiering och programplanering för kulturellt samarbete ( kultur 2000-programmet ) c5-0327 / 1999 - 1998 / 0169 ( cod ) ) .
fru talman ! jag tror egentligen att vi inte hade behövt tala mer om det , ty vi har redan sagt allting under den senaste debatten .
tyvärr har ju ingenting ändrats i fråga om det faktum att rådet alltid talar om kultur , men inte ger ut några pengar för kultur .
vi har en känsla av , och är egentligen övertygade om , att medlemsstaterna skulle uppskatta om de kunde stryka det som de 1992 skrev in i maastrichtfördraget .
ty ingen vill egentligen verkligen ge ut pengar för kultur .
tyvärr är det så . det måste vi konstatera .
jag vill tacka föredraganden , som verkligen oförtröttat har arbetat med detta omfattande ärende , naturligtvis i samarbete med kommissionären .
vi måste nog notera att vi egentligen har uppnått vårt mål beträffande innehållet , men naturligtvis inte beträffande finanserna .
i en sådan förlikning , där man å ena sidan verkligen måste uppnå enhällighet , känner man sig maktlös .
det är egentligen inte någon rättvis basar !
det finns alltid människor där som kan avvisa allting , och å andra sidan står vi och tigger om lite mer för kulturen .
det är egentligen vanhedrande , det som vi gör där !
det är en förskräcklig arabisk basar , med ojämna förutsättningar .
det gläder oss ändå att detta program har blivit sådant som vi önskade .
det motsvarar det som medborgarna förväntar sig av oss .
vi stöder små och medelstora arrangemang , inte de stora arrangemangen , vi gör tillgången till det enklare för den enskilde medborgaren och även de mindre aktörerna ; jag tror att det faktum att kulturen i dag ju tillsammans med utbildning och ungdom befinner sig i en kommissionärs hand , också borgar för att det skapas mer synergi mellan dessa tre program , som ju är utpräglade program för medborgarna i europeiska unionen .
om man tar alla pengar och åstadkommer synergieffekter , då kan man var litet tillfreds , men också bara litet grand .
jag önskar att vi med dessa mindre summor uppnår många effekter .
fru talman ! jag håller med om de stora ord som fick inleda föredragandens anförande , men jag måste få tillägga att jag under förlikningen har blivit lite besviken på rådet .
å ena sidan vägrade man fortfarande att acceptera begreppet &quot; europeisk kulturpolitik &quot; och liknande begrepp , bland annat genom att förringa det som står i fördragen , och man har endast definierat begreppet &quot; kultur 2000 &quot; som ett instrument för ett kulturellt samarbete , och mer än så blir det inte .
å andra sidan har man visat sig helt omedgörlig beträffande den finansiering som parlamentet har begärt , som gällde en minimifinansiering .
nåja , det vore orättvist att påstå att det sista rörde rådets fjorton medlemmar , för det var bara en , nederländerna , som i första hand visade sig omedgörlig .
det har än en gång visat sig att en förlikning är oförenlig med kravet på enhällighet i rådet .
ett sådant krav gör i princip en förlikning omöjlig och inverkar dessutom på den parlamentariska institutionens värdighet .
fru talman , dessa överväganden får emellertid inte dölja det faktum att denna text som i sin helhet kommer att bli föremål för omröstning i morgon , och som vi socialister kommer att rösta för , kommer att innebära igångsättandet av ett av europeiska unionens viktigaste program .
genom att agera på det kulturella området , skapar vi europas själ , inte minst i det här fallet med de fantastiska gemenskapsprogram som utgör &quot; kultur 2000 &quot; .
de senaste åren har dessa blivit de mest accepterade programmen bland de mest dynamiska och yngsta medborgarna i europeiska unionen .
slutligen vill jag nämna det starka intryck som föredragande graca moura som individ har gjort på mig : hans kunskap , hans eftertanke , hans intellektuella nivå visar , anser jag , att han är den bästa föredraganden som detta betänkande hade kunnat få .
till sist vill jag gratulera kommissionär reding , vice talman imbeni samt gargani , ordförande i utskottet för kultur , ungdomsfrågor , utbildning , medier och idrott , för den bestämda och kloka hållning som de , var och en i sin roll , har intagit under hela förlikningsprocessen .
fru talman , fru kommissionär , herr föredragande ! jag skulle vilja börja med att tacka graça moura så hjärtligt för hans fantastiska insats under behandlingen av programmet kultur 2000 .
det har redan sagts och vi har diskuterat det flera gånger , kultur är naturligtvis otroligt viktigt som ett självständigt område , det vill jag betona igen , men också som ett utmärkt instrument för att vidarebefordra den europeiska tanken och kulturen är mycket viktig för medborgarna .
det får vi absolut inte glömma bort .
det europeiska stimulans som ges ut genom det här programmet medför otroligt mycket , särskilt för små språkområden som t.ex. nederländerna där det inte endast gäller nationella möjligheter men de behöver också stödjas , framförallt genom språket .
i dag har vi kommit fram till slutet av en lång resa .
jag skulle ändå helt kort vilja , precis som andra gjort , gå in på det otydliga och främst ovälkomna förfarandet .
medbeslutande och enhällighet är som en orm som biter sig själv i svansen .
det finns inte mycket att förhandla om i fall en av parterna på förhand säger : vi kan prata om allt men budgeten står fast .
nu har , och det vill jag ändå också säga när det gäller nederländerna , förhandlingarna om det redan ägt rum i ett tidigare skede .
resultatet är 30 procents tillväxt , så vi är inte helt olyckliga över resultatet .
det är naturligtvis alltid bättre , och det skall jag alltid yrka för , att anslå mer pengar och även något snabbare . ändå så tror jag att det här programmet erbjuder goda chanser för flera olika program .
jag skulle vilja betona att kultur inte enbart får stöd från den här fonden .
kultur består inte enbart av kultur utan även av många andra områden .
i strukturfonderna finns också mycket pengar tillgängliga för kultur och det måste vi ju också ta i gott beaktande .
lyckligtvis är jag ledamot i utskottet för regionalpolitik .
jag skall alltså själv se till att det också sker i stor utsträckning .
jag tror att vi även tagit ställning för att instämma i att budgeten är tillräckligt omfattande , om det inte går igenom så är det ju ändå dåligt för medborgaren .
i det avseendet har jag också alltid stöttat föredraganden .
jag tycker dock att det , och det säger han också alltid , vid den kommande regeringskonferensen behöver göras en ändring i medbeslutandeförfarandet , då behövs ingen enhällighet .
vi är mycket positiva över de många förbättringar som skett . inga megaprojekt längre , utrymme för kulturella nätverk , god uppmärksamhet för läsfrämjande åtgärder , översättning , översättarhus , mycket viktigt för de mindre språkområdena .
jag vill verkligen lyckönska föredraganden och även reding till kultur 2000 .
det enda som återstår för mig att säga är : nu sätter vi igång .
fru talman ! de kolleger som har talat före mig har sagt det mesta , och jag tror att det finns en samstämmighet bland grupperna i europaparlamentet liksom bland alla oss i utskottet för kultur , ungdomsfrågor , utbildning , medier och idrott .
även jag skall säga att det är med ett mycket tungt hjärta som jag kommer att rösta för detta gemensamma förslag till rådets och europaparlamentets beslut .
inte på grund av att våra företrädare , vår föredragande och ordföranden gargani , inte har uträttat ett enastående arbete - det har lagt ned enormt mycket arbete - , inte på grund av att jag har några stora invändningar mot den ståndpunkt som kommissionär reding har vidhållit - jag tycker att hon inom de ramar som hon hade vidhöll en mycket positiv ståndpunkt - , utan på grund av rådets negativa och oacceptabla inställning .
det är en skam !
denna siffra , 167 miljoner euro för så många år , är en skam för europeiska unionen !
när vi bokstavligen tvingas att kväva teatergrupper , unga musiker , innovativa verksamheter inom konst och litteratur , att kväva dem och hålla god min och ge femtioelva avslag , med resultatet att de uppfattar europa som någonting främmande , någonting motsträvigt , någonting negativt och någonting fientligt i sina ansträngningar att skapa kultur , ansträngningar som europeiska unionen måste stödja - för vår väg är inte bara euron , inte heller bara utvidgningen eller egoistiska geostrategiska hänsyn ; den är att ge en kulturell blomstring till den europeisk integrering - , är denna utgång beklaglig .
och så länge som vi har kvar enhälligheten och så länge som en regering , som nederländernas regering i går , kan fastställa de där 167 miljonerna med ett ultimatum och så länge som en regering med haider i övermorgon kan tala om för oss vilka kulturella verksamheter vi skall ägna oss åt , kommer vi inte att komma framåt .
därför är det mycket viktigt för regeringskonferensen att det fattas viktiga beslut och att det kommer till stånd en ändring , så att europaparlamentets ansträngningar att få till stånd en viktig kulturell blomstring inom det europeiska området befrias från enskilda regeringarnas tvångströjor .
fru talman ! jag delar helt de värderingar som har framförts av föredraganden och jag vill också tacka ordföranden för utskottet för kultur , gargani , för det berömvärda arbete han utfört under en medlingsprocess som även varit ganska komplicerad .
utan tvekan finns det behov av att förenkla och förstärka tidigare program men alla hoppades att programmet kultur 2000 skulle kunna bidra till att till exempel främja varje kultursektors särart , och även - eller framför allt , bör man kanske säga - de sektorer som inte är så kända .
vi hoppas att detta skall inträffa , åtminstone när det gäller finansieringen .
vi tror mycket på värdet av kulturella handlingar , även när det gäller bidragen till ett folks sociala och ekonomiska tillväxt .
och europa kan fullt ut konkurrera med resten av världen genom att till fullo återupptäcka sina rötter , genom att förverkliga det gemensamma kulturella nätverket , genom att utnyttja och återge värdigheten åt de kulturella och språkliga öar som hittills varit mindre kända .
när det gäller den stora pedagogiska uppgift som europeiska unionen står inför i samband med den kulturella dimensionen , är finansieringen en av de tydligaste begränsningarna när det gäller programmet - det har vi fått höra flera gånger - och något som pekar på att man inte har helt förstått - åtminstone gäller det rådet , men sannerligen inte kommissionären - betydelsen av denna kulturella uppgift : detta visar även dokumentet som prioriterar de ekonomiska faktorerna framför den sociala integrationen .
en allsidig tillväxt av europeiska unionen och medvetenhet om vad det innebär att vara europeiska medborgare : det är därför vi anser att projektet kultur 2000 , även när det gäller finansieringen , skulle kunna lämna viktiga bidrag till detta stora gemensamma mål .
fru talman ! jag vill öka kvällens enhällighet och säga att jag stöder godkännandet av kultur 2000 och framför mina tack till föredragande , graca moura , som efterträdde vår förra kollega nana mouskouri .
båda har gjort ett förstklassigt arbete .
vid sidan av den debatt vi hade tidigare i dag kanske kultur inte verkar vara så viktig men den är det och vi måste vara varsamma i europaparlamentet så att brådskande frågor inte går före vad som är viktigt .
varför anser jag att kultur är viktig ?
jo , i enkla ekonomiska termer främjar europeisk kultur verkligt välstånd .
var skulle europas turistindustri befinna sig utan rikedomen i vår kultur ?
men viktigare än det , kulturaktiviteter är det som gör människosläktet civiliserat .
kulturen är grunden för vår tro på demokrati och ett icke kulturellt samhälle kan inte upprätthålla tolerans och frihet och demokrati .
kulturell mångfald är viktig och den är hotad .
men hotet kommer inte från europa .
många människor i mitt land säger att de uppfattar att brittisk kultur hotas exempelvis från portugal , tyskland , finland , för guds skull .
vi dricker ju portvin och vi tycker om tyskt öl och vi använder till och med finsk bastu men det är inte från europa som kulturen hotas .
vad jag verkligen ser i hela europa är folk som dricker coca cola , som äter hamburgare , bär baseballmössor , tittar på hollywoodfilmer och ofta gör allt detta samtidigt .
jag tror inte att protektionism och reglering är rätt metod för att försvara europas kultur , men jag tror att vi ska ge en hjälpande hand när vi har möjlighet .
det är vad kultur 2000 handlar om .
så jag säger till ministerrådet : utvärdera verkligen ständigt detta program .
gör vi tillräckligt mycket ?
och jag säger till fru reding , tack för det stöd och den hjälp ni har gett hittills , fortsätt göra ett bra jobb , vi står på er sida .
fru talman ! även jag vill varmt tacka föredraganden graça moura och kommissionsledamoten reding för deras ansträngningar för att åstadkomma detta program .
kultur 2000-programmet fick ju sin slutgiltiga form i slutet av förra året genom förlikningen mellan parlamentet och rådet .
slutresultatet kan anses vara rimligt med tanke på att det krävdes ett enhälligt beslut i rådet för att godkänna programmet .
det är önskvärt att man vid den kommande regeringskonferensen kommer fram till att införa beslut med kvalificerad majoritet även inom kulturens område .
det är verkligen besynnerligt att lagstiftning där man tillämpar medbeslutandeförfarandet förutsätter enhällighet i rådet .
det kulturella ramprogrammet ersätter de nuvarande programmen kalejdoskop , ariane och rafael .
när man börjar genomföra programmet hoppas jag speciellt att möjligheterna för litteraturen och översättningen av böcker kan utnyttjas fullt ut .
jag tror och hoppas att litteraturen bibehåller sin ställning trots den nya teknikens framfart .
vi behöver den fördjupning som litteraturen erbjuder mitt i all kortsiktighet och ytlighet .
litteraturen har likaså en stor betydelse när det gäller att förmedla vårt kulturarv , att öka kännedomen om varandra samt att omhulda den språkliga rikedomen och mångfalden .
i detta sammanhang är det speciellt angenämt att konstatera att eu : s ordförandeland strax efter att sokrates- och kultur 2000-programmet startats kommer att anordna ett möte där man skall dryfta bibliotekens ställning .
jag hoppas att detta möte också skall uppmuntra kommissionen till att på ett aktivt sätt beakta biblioteken i informationssamhällets femte ramprogram .
fru talman , fru kommissionär , herr föredragande , mina damer och herrar ! någonstans sluts kretsen med dagens föredragningslista .
vi har i dag talat mycket om europa som en värdegemenskap , om tolerans , mänsklig värdighet , mänskliga rättigheter , ett positivt förhållande till utvidgningsprocessen , öppenhet och respekt för varandra .
ungdoms- , utbildnings- och kulturpolitik är viktiga verktyg när man skall skapa dessa värden , skapa förtroende hos medborgarna i europeiska unionen och skapa trovärdighet för europeiska unionen gentemot medborgarna .
de finansiella medel som av rådet medgivits för kulturprogrammet står i ett slående motsatsförhållande till betydelsen av kultur- och utbildningspolitiken samt detta program för europeiska unionens mål .
kulturell verksamhet skapar identitet .
kulturell verksamhet är ett uttryck för individualitet och den egna personligheten , den skapar kontakt och kommunicerar .
vi vill ha ett brokigt europa .
vi vill ha ett europa enligt principen mångfald inom enheten .
vi vill att människorna skall lära sig förstå och uppskatta skillnaderna .
av den anledningen har vi uttalat oss för en uppdelning av budgeten respektive anslag till de olika typerna av åtgärder .
av den anledningen har vi avvisat den starka koncentrationen till stora nätverk och nätstrukturer , eftersom vi vill främja de små och medelstora enheterna , den individuella verksamheten , eftersom vi vill låta tusen blommor blomma .
jag vill stödja de föregående talarna .
det är en motsägelse - enhällighetsprincip , medbeslutandeförfarande och förlikningskommitté - om vi vill stärka kulturpolitikens principer för ett europeiskt medvetande och inte vill fortsätta att försvaga dem .
fru talman , mina damer och herrar ! som vi har hört , har alla våra grupper en gemensam politisk fiende , och det är rådet .
utskottets för kultur beslut hamnar ju inte av en tillfällighet alltid i ett förlikningsförfarande , ty det är alltid något medlemsland i rådet som tar kulturen till gisslan för andra intressen .
så visar sig enhällighetsprincipen vara ett första klassens blockadinstrument .
i nästan två år har man brottats för att uppnå en genomförbar kompromiss , innan europaparlamentet nu äntligen kan ge grönt ljus .
inte ens det faktum att de föregående programmen kaleidoskop , ariane och rafael löpte ut kunde beveka rådet .
det krävdes ett pilotprogram för att överbrygga detta .
det har än en gång tydliggjort svagheterna i europeiska unionens kulturpolitiska åtgärder .
den politiska kampen om anslagsfördelningen och programutformningen står inte i någon proportion till volymen på stöden .
av 410 framställningar år 1999 kunde bara 55 projekt med en mager totalvolym om 6,07 miljoner euro beaktas .
beträffande föreliggande program var rådet inte berett att komma parlamentet till mötes med en enda euro !
alltså stannar vi kvar på blygsamma 167 miljoner till år 2004 .
det motsvarar utgifterna för ett enda medelstort tyskt operahus under samma period , medan denna summa här i europa är avsedd för 29 länder i över 5 år .
det är ett krasst missförhållande !
alltså måste vi då vredgat finna oss till rätta med att vi åtminstone i fråga om innehållet har fått igenom en del .
det har ju också redan lyckligtvis skildrats .
hoppet kvarstår att det en dag kommer att bli möjligt att förmå rådet att ändra inställning .
kanske kommer man ju också att begripa att europeiska unionens kulturella aktiviteter inte utgör någon fara , utan en möjlighet !
kulturellt samarbete - även detta har skildrats - bidrar sannerligen till att ge en identitet , mycket mer än alla viktiga transportdirektiv .
att man främjar kulturen bemöts med allmän acceptans , vilket man sannerligen inte kan påstå om alla politiska beslut .
vad är det alltså , frågar jag er , som rådet är ängsligt för ?
fru talman ! den som , i likhet med mig , har äran att vara ordförande för kulturutskottet kan inte annat än instämma i det som har sagts av diverse kolleger och jag kan inte låta bli att gratulera föredraganden och kommissionären , fru reding , med vilken föredraganden har arbetet och som , även i förlikningen , har haft svåra stunder , har kämpat mot rådet , det har vi fått höra av alla .
jag har kunnat konstatera hur starkt man har bekräftat principen om kulturens nödvändighet när det gäller det europeiska konstruktionsarbetet men med små möjligheter att tillfredsställa alla de krav som kommer från europas olika stater .
låt mig bara understryka mitt personliga beklagande över att man i slutändan inte har lyckats godkänna en revideringsklausul .
vi har , det är sant , fru redings villighet och långsiktiga mål , reding som har engagerat sig personligen för att ta upp frågan på nytt , för att göra en heltäckande utvärdering om något år , och därmed få till stånd en ny situation .
de olika kulturprogram - kaleidoskop , ariane , rafael - som har startats under de år som gått ersätts nu av ett enda program , kultur 2000 , där - detta vill jag gärna understryka - föredraganden stigmatiserat en åsikt som borde få europaparlamentet att tänka efter - vilket någon redan påpekat under eftermiddagen i dag - men som alltid understryker den stora betydelsen av att vara del av en stor gemenskap där kulturen är ett demokratiskt fenomen .
detta är ingen tom retorik , utan snarare en ny typ av liberalism som förenar de europeiska staterna och som är en utmaning för europaparlamentet och kommissionen .
vi har enats i den här frågan och det resultat som vi i dag har uppnått , trots den bristfälliga finansieringen , tror jag kan göra så att denna strategi och denna möjlighet för europa verkligen får en bred lansering , en strategi som kommer att bli avgörande för såväl ekonomin som utvecklingen : med andra ord kulturen , ett institutionellt och organisatoriskt faktum som en förutsättning för den ekonomiska utvecklingen , och inte tvärtom , som europa av tradition tyvärr har haft för ovana att se det under de år som gått .
i första hand handlar det om människan , i första hand handlar det om kulturen , och den kulturen kan avgöra den ekonomiska utvecklingen .
låt oss begrunda detta resultat , låt oss vara glada och låt oss ge oss själva stor frihet att utforma en användbar strategi .
fru talman ! får jag först och främst tacka herr graça moura för att ha vävt sin väg genom de ganska hårda vävnader och trådar som denna förlikningsvävnad bestod av .
det förefaller mig när vi inledde förliknings- förfarandet för kultur 2000 att det är helt passande att ha en poet att leda oss i vår strävan .
då dessa förlikningar inte utvecklas i helt rak kurs måste vi på nytt tacka vice talman imbeni för hans föredömliga förhandlingsskicklighet på det invecklade området för att se till att kulturanslag sprids ut på ett klokt sätt och ges till oss i vår gemenskap .
jag tycker att den huvudfråga som detta parlament , kommissionen och rådet står inför verkar vara : vad är europa ?
vad betyder europa och vad ger europa oss utöver parametrarna för våra nationella gränser ?
europa är dess folk , dess historia och nu dess gemenskap . skälet till varför kultur 2000 är så viktig för oss är emellertid detta : jag skall slå vad om det när vi ställer frågan - &apos; vad är europa ?
vi svarar med att säga : &quot; det är vår konst , det är vår litteratur och det är vårt arv . &quot;
det är vad kultur 2000 står för . detta program står för möjligheten att bibehålla en europeisk identitet på 2000-talet , en identitet som saknar ekon av splittring , av krig , av fattigdom , av möjligheter , av fattigdom i verkligheten .
och mer än detta - och detta är mer vardagligt , fru talman , innebär det att vi har förmåga att lära från tidigare politiska initiativ genom att tillämpa dem i nya program som är innehållsrika , som täcker flera områden och som är till nytta för våra kreativa industrier i den utsträckning som de nu behöver .
det främjar rörlighet och öppnar dörrar till kultur för de socialt missgynnade och utslagna .
det enda jag beklagar är att vi inte har tillräckligt med pengar för att stödja detta program i överensstämmelse med våra förhoppningar och så att vi kan säkerställa att vi kommer att kunna nå ända fram .
( fr ) fru talman , mina damer och herrar ! vi har nu kommit till slutet på en lång väg .
efter förlikningsetappen kan våra institutioner numera formellt anta det nya ramprogrammet &quot; kultur 2000 &quot; .
vi förfogar då över ett instrument som gör det fullständigt möjligt att under de fem kommande åren utveckla en tydlig och väl strukturerad och , det är jag säger på , lönsam åtgärd , till förmån för kultursektorn .
det är med tillfredsställelse jag i dag här välkomnar denna happy end och jag tackar er .
jag tackar alla dem som här i parlamentet arbetat för att en bra avslutning på förlikningen kunnat bli möjlig .
jag vill uttrycka mitt tack särskilt till utskottet för kultur , ungdomsfrågor , utbildning , medier och idrott och bl.a. dess föredragande graça moura , dess ordförande gargani , till europaparlamentets delegation och de ansvariga för de politiska grupperna , till förlikningskommittén och dess ordförande imbeni .
alla har bidragit konstruktivt , rättvist och beslutsamt .
under hela denna förhandling har de varit till stor hjälp och det måste sägas att den svåra , ibland smärtsamma , förhandlingen ändå genomförts på rekordtid .
vi har nu ett ramprogram , det första i detta slag för kultursektorn , och detta program gör det möjligt för oss att planera våra åtgärder ur en ny synvinkel och arbeta till förmån för kulturen på ett mer globalt , men också mer komplett och mer fördjupat sätt .
jag gläds med er åt dessa tillfredsställande resultat som måste göra det möjligt för oss att , trots en budgetsituation som inte ligger i nivå med våra ambitioner , se framtiden an på ett mycket positivt sätt , och jag skulle vilja ta upp det som ordförande gargani sade : kommissionen har gjort ett uttalande beträffande utvärderingen efter halva tiden .
den har förklarat att i samband med den rapport den måste utarbeta i enlighet med artikel 7 i beslutet från parlamentet och rådet kommer den att genomföra utvärderingen av programmets resultat , och denna utvärdering kommer även att gälla de ekonomiska resurserna inom ramen för gemenskapens budgetplan .
vid behov kommer rapporten att innehålla ett förslag till ändring av beslutet och allt detta före den 30 juni 2002 .
mina damer och herrar , kära parlamentsledamöter ! det är ett formellt åtagande , inte bara en mening på ett papper .
allt detta måste leda oss till att stärka våra åtgärder till förmån för att lyfta fram ett gemensamt kulturområde , inom vilket våra kulturer kan utvecklas ytterligare i alla sina specifika karaktärer , all sin mångfald , men de kan också berikas ömsesidigt och övriga europeiska medborgare kan delta fullt ut .
det är också tack vare parlamentet som vill att fler små åtgärder skall genomföras nära medborgarnas rötter snarare än stora spektakulära åtgärder .
detta kommer att leda till att vi gör programmet &quot; kultur 2000 &quot; till ett program för medborgarna .
detta ökade deltagande från medborgarnas sida , som jag verkligen hoppas på , vill jag skall vara så brett och fruktbart som möjligt och jag förbinder mig att verka för att det blir en nåbar verklighet under de fem år som omfattas av programmet .
jag vet att ni parlamentariker , i era regioner , i era länder , kommer att verka tillsammans med deltagarna i programmen för att alla dessa små blommor , som en kollega sade , skall bli en stor mångfärgad matta .
jag skulle vilja att detta program blir en nåbar verklighet och att kulturen för våra medborgare utgör inte bara en berikande faktor , såväl på det personliga som det sociala och ekonomiska planet , utan även en rättighet som det handlar om att bekräfta , liksom ett tecken på en återfunnen sällskaplighet inom unionen .
det är vad vårt europeiska program &quot; kultur 2000 &quot; tillför .
det är inte någon konkurrent till den kulturpolitik som bedrivs i de olika medlemsstaterna .
den är nödvändig och jag skulle vilja se den utvecklas ytterligare .
det är helt enkelt ett tillägg , ett komplement , ett byggande av en bro mellan de olika kulturerna i våra olika länder .
att utvidga och berika de europeiska medborgarnas deltagande i kulturen förefaller mig alltså vara en grundläggande uppgift som motiverar våra ansträngningar och hur vi bör bedöma framgången med vår åtgärd och med vår union .
flera parlamentariker har med rätta tagit upp det : om en union enbart består av ekonomi är den dödfödd .
men om den består av kultur , om den består av civilisation , om den består av deltagande kommer den att bli levande .
det är denna grund , mina damer och herrar , som jag har för avsikt att utveckla och jag kommer särskilt att ta hänsyn till följande inriktningar : för det första erbjuda möjligheter av innovativ karaktär för våra kreatörer så att deras talanger får det stöd de förtjänar i vårt program .
för det andra uppmuntra utbyte , rörlighet , utbildning inom kultursektorn .
för det tredje främja samarbete mellan kulturarbetare .
för det fjärde utöka allmänheten genom att bl.a. göra större plats för ungdomarna , och för det femte bevara och göra det gemensamma kulturarvet av europeisk betydelse mer känt , liksom de europeiska folkens historia .
det nya programmet blir , genom sin struktur , sin organisation grundad på öppenhet , effektivitet och balans , det är jag säker på , ett instrument med lika hög prestanda som det blir grundläggande för våra åtgärder .
fru talman ! jag upprepar mitt tack till parlamentet för dess stöd och för att ännu en gång ha visat på den betydelse det fäster vid kulturen i unionssammanhang .
jag är övertygad om att parlamentet inte kommer att bli besviket för att ha beviljat oss sitt stöd och jag förbinder mig att personligen successivt informera parlamentet om olika etapper i genomförandet av våra åtgärder , våra medborgares åtgärder , som jag hoppas skall bli stora åtgärder för unionens framtid .
jag tror att vi kan tacka vår föredragande ännu en gång .
( sammanträdet avslutades kl. 21.55 )
uttjänta fordon
nästa punkt på föredragningslistan är andrabehandlingsrekommendation ( a5-0006 / 00 ) från utskottet för miljö , folkhälsa och konsumentfrågor om rådets gemensamma ståndpunkt ( 8095 / 1 / 1999 - c5-0180 / 1999 - 1997 / 0194 ( cod ) ) inför antagandet av europaparlamentets och rådets direktiv om uttjänta fordon ( föredragande karl heinz florenz ) .
herr talman , ärade damer och herrar , kära kolleger ! årligen skrotas nio miljoner bilar i europa .
trots det faktum att dessa nio miljoner bilar inte längre kan köras har de den egenskapen att man handlar med dessa även mindre legalt även över gränserna , inte bara över gemenskapens inre gränser utan även över gränser som ligger utanför unionen .
därför är det principiellt riktigt att europeiska unionen upprättar allmänna spelregler för hur dessa nio miljoner fordon per år skall återvinnas och tas om hand .
direktivet har enligt oss ett par svagheter som vi gärna vill rätta till här i kammaren genom ett direktiv som då verkligen blir framtidsinriktat .
därför finns det en mängd ändringsförslag .
jag personligen anser att man genom direktivets tillämpningsområde skjuter över målet .
jag anser det inte nödvändigt att veteranbilar skall utgöra en del av direktivet .
jag tycker heller inte att motorcyklar bör omfattas av direktivet , eftersom återanvändningen i fråga om motorcyklar är en så särskild kulturform att det inte behövs några europeiska direktiv för detta .
inte heller för specialfordon eftersträvar jag nödvändigtvis höga återanvändningsnivåer .
min önskan är den att specialfordon såsom ambulanser skall nå höga räddningsnivåer .
det är mitt huvudsakliga bekymmer på det området .
återvinningskraven på hur avfall från bilar skall hanteras i europa föreskrivs efter mitt förmenande på ett bra sätt i direktivet .
här kan det få stanna vid det som kommissionen har föreslagit .
medlemsstaterna sörjer för att det finns motsvarande insamlingsanläggning där man tappar ur bilarna , tar hand om exempelvis över 32 miljoner spillolja , tömmer dem på bromsvätska etc.
en viktig komponent i direktivet är frågan : vad vi skall göra med de gamla bildelarna ?
vad gör vi med de skrotade produkterna ?
man får inte blunda för att det kvantifierade målet är en viktig punkt när det gäller recycling ( återvinning ) och återanvändning ( recovering ) och vad det nu är , men det är inte den enda punkten .
för vi skall inte glömma : under en bils livscykel faller 80 procent av miljöbelastningen på körningen , 1 procent på sluthanteringen och 19 procent på tillverkningen av bilen .
kvantifierade målsättningar är sålunda inte den enda parametern vid frågan om miljökonsekvenserna , utan en av många .
jag är naturligtvis av den uppfattningen att vi behöver rigorösa mål .
men kvoterna får inte bli ett självändamål , utan vi måste inse att helhetssynen på hur bilen belastar miljön är viktig .
jag ser mycket hellre att vi kommer bort från en bil som i dag väger 1 400 kilo , som körs i genomsnitt i 200 000 km , till en bil som i framtiden väger endast 1 000 kilo och också körs i 200 000 km .
trots allt skulle det då transporteras 400 kilo gånger 200 000 km mindre .
detta är det sanna miljöpolitiska framsteget , för det leder till en kraftig minskning av koldioxid och detta är , om jag har förstått kyotoprotokollet rätt , den viktiga beståndsdelen .
därför tror vi att fordon som i framtiden på ett imponerande och påvisbart sätt använder sig av lättviktsmetoder producerar mindre koldioxid och ges speciella preferenser i förbränningskvoten .
detta skall inte den enskilda medlemsstaten besluta om , utan det är ni , fru kommissionär , som tillsammans med er stab skall besluta om huruvida dessa lättviktsfordon - många talar även om 3-liter-bilar - skall erhålla speciella preferenser .
vi är av den uppfattningen att det är riktigt .
låt mig säga något om kostnaderna .
vissa säger att tillverkarna borde få bära hela kostnaden - det skulle vara riktigt och mycket konsumentvänligt .
detta kan man ifrågasätta mycket starkt , för tillverkarna kommer att lägga över alla kostnader på konsumenterna och tillägna sig ett återvinningsmonopol som borde vara statligt .
jag kan bara varna er för att rösta för detta .
det finns ändringsförslag som går ut på att kostnaderna skall delas , hälften åt tillverkarna och den andra hälften åt nybilsköparna .
ur en sådan pool , ett sådant system , hur ni nu än föreställer er detta , kan man då från och med 2006 återta alla fordon i bilparken utan kostnad för den sista ägaren .
detta är också min grupps uttryckliga önskan .
vårt förslag om delning av kostnaderna har en alldeles avgörande fördel , nämligen att vi slipper bli domstolskandidat så snart vi har antagit direktivet .
för den återverkan som bilindustrin så listigt betalar tillbaka med är ett allvarligt problem som vi rimligen måste ta hänsyn till .
därför föreslår jag att kostnaderna delas av den första ägaren och tillverkaren .
förbud mot vissa material - naturligtvis behöver vi förbud mot vissa material .
det finns farliga komponenter i bilen , dessa måste på sikt förbjudas .
till det behöver vi ett instrument för påtryckningar .
kommissionen har lagt fram några förslag som var för stränga , och vi har tagit fram alternativ till dessa .
det finns en mängd bra ändringsförslag .
parlamentet har fått större befogenheter . så låt oss utnyttja dessa !
låt oss vara modiga nog att lägga fram och utveckla ett direktiv som pekar in i framtiden .
ett direktiv som utvecklas endast för direktivens egen skull vore inte värdigt kammaren .
herr talman , fru kommissionär , kära kolleger ! när man ser de flygblad som har delats ut under de senaste veckorna så tror man att det är en möjlig miljökatastrof eller den europeiska bilindustrins död vi diskuterar här. inte något av detta stämmer .
vi måste se med nyktra ögon på att direktivet som ligger framför oss på bordet är ett bra direktiv .
det innebär miljömässiga framsteg för europa , och vi kan vara stolta om vi kan få till stånd och förankra direktivet i lag .
förvisso , det finns en punkt som vi är oense om .
med tanke på direktivets dimensioner är det måhända en liten punkt , men det är detta oenigheterna handlar om .
det gäller frågan om kostnaderna för återvinningen .
här skiljer vi oss i väsentliga delar från diskussionen i rådet förra året . där drogs nämligen kostnadsbefrielsen för sista ägaren och frågan om finansieringen över en kam , och kostnadsbefrielsen för sista ägaren ifrågasattes .
vi här i kammaren fattade entydigt beslut i februari förra året - och detta stöder vi , just vi socialdemokrater - kostnadsbefrielsen för sista ägaren är för oss odiskutabel !
men vem betalar för de fordon som skall skrotas och tas om hand ?
för oss är det självklart att tillverkaren skall göra detta vad gäller nya bilar , därför att detta också är ett incitament för tillverkaren att ta fram och tillverka återvinningsvänliga bilar .
men vad händer med fordonen som rullar på gatorna ?
ett exempel : firman rover i storbritannien skulle , om man blev ansvarig för alla uttjänta fordon , bli ansvarig för 5,8 miljoner bilar i europeiska unionen och omgående tvingas öronmärka 250 miljoner euro för att spara ihop till återvinningskostnaderna , medan en tillverkare av liknande bilar från korea behöver lägga undan ett peanuts-belopp - som en företrädare för deutsche bank en gång uttryckte det .
här finns en snedvridning av konkurrensen som inte har med miljöskyddet att göra utan enbart inverkar på investeringsförmågan , och på arbeten för de människor som bygger bilar här i europa .
i så måtto föreslår jag att en fond för de gamla fordonen bildas , ur vilken återvinningskostnaderna för de uttjänta fordonen sedan betalas så att principen om kostnadsbefrielse säkras .
jag kan förstå att kolleger från länder utan biltillverkning säger ja , tillverkarna skall betala alltihop , och problemet med snedvridningen av konkurrensen genom öronmärkta reserver intresserar oss inte !
men jag ber dessa kolleger visa solidaritet med de drygt två miljoner människor som tillverkar bilar i europa , som på så sätt finansierar sina liv , så att dessa arbetsplatser kan garanteras även i framtiden .
jag är för stränga miljökrav , det vet ni från auto / oil-programmet och diskussionen om gränsvärdena för avgaser . men jag anser att kraven måste vara lika för alla !
herr talman , herr kommissionär , kolleger ! jag tror att vi behöver detta direktiv .
för det första eftersom det innehåller en tydlig beskrivning av miljömålsättningarna .
för det andra eftersom detta direktiv kan stimulera återanvändning , och det är viktigt .
för det tredje finns det ett tydligt tillvägagångssätt för att motverka föroreningen från tunga metaller .
det är också en viktig punkt .
direktivet ger en europeisk ram , bland annat också för medlemsstater som redan har ett system och som vill fortsätta att arbeta med det systemet .
vi måste således i första hand bibehålla procentandelarna i fråga om återvinning , för därigenom uppmuntrar man naturligtvis teknisk förnyelse och olika sätt att hitta en lösning för material som vi ännu inte riktigt vet vad vi skall göra med .
för det andra måste vi låta de omständigheter som står i den gemensamma ståndpunkten vara oförändrade .
så från och med år 2006 gäller kostnadsfri inlämning för alla bilar , kostnadsfri för den sista ägaren .
det är naturligtvis helt klart en mycket viktig punkt . den får vi inte tumma på .
är detta en för stor börda ?
det finns dock en sak som vi inte får glömma bort .
direktivet handlar om fullständiga bilar , alltså bilar där inga viktiga delar saknas .
enligt experterna är det inte många av dessa fullständiga bilar som är värdelösa .
för återvinning , återanvändning av delar , det är en sektor som inte nödvändigtvis är förlustbringande .
tvärtom , det finns för närvarande ett stort antal företag som lever av detta och som därigenom utan problem kan förtjäna sitt levebröd .
detta direktiv stimulerar hela denna sektor .
det handlar om en sektor som utgörs av små och medelstora företag .
eftersom transportkostnaderna i detta fall ligger på en hög nivå måste det också bli fråga om ett starkt decentraliserat system , för att flytta ett vrak mer än 100 kilometer är inte någon lönsam verksamhet .
jag tycker att det är en bra idé att detta direktiv inte skall gälla för historiska bilar , och jag anser att det måste vi lägga till .
så enligt min uppfattning bör veteranbilar befrias från detta .
det är också bra att vi tydligt lägger ansvaret hos producenten .
det är en grundläggande princip och den måste vi hålla fast vid .
han är ansvarig för konstruktionen . han kan således göra en mycket stor insats för miljön i samband med denna konstruktion .
vi måste också hålla fast vid att kostnaderna skall bäras av producenten , helt eller till övervägande delen , vilket står i den gemensamma ståndpunkten .
jag anser att det är en balanserad princip som inte utesluter några andra saker .
min uppfattning är att vi måste behålla denna .
därför kommer vår grupp att stå kvar så nära den ursprungliga gemensamma ståndpunkten som möjligt och inte förändra denna ståndpunkt på de väsentliga punkterna .
för vi vet naturligtvis allesammans att det var mycket mödosamt att få till stånd denna ståndpunkt i rådet , att det var en svår balansövning att uppnå denna gemensamma ståndpunkt .
vi får , enligt min uppfattning , från vår sida inte sätta denna gemensamma ståndpunkt i fara , för detta är ett direktiv som vi absolut behöver av miljöskäl .
jag uppmanar er att stödja denna gemensamma ståndpunkt .
vår grupp kommer i vilket fall att göra detta i så stor utsträckning som möjligt av miljöskäl eftersom vi har detta direktiv och eftersom det är ett balanserat direktiv som innehåller en mängd saker , en mängd invändningar , till exempel i fråga om kostnadsfördelningen .
herr talman , kolleger ! i dag har vi ett viktigt beslut att fatta .
stöder europaparlamentet den ekologiska principen om producentansvar , det vill säga att fordonstillverkarna har ansvaret för bilar när de har blivit bilvrak ?
nej , säger kristdemokraterna i ändringsförslag 38 : fordonstillverkare och bilister skall dela kostnaderna lika .
i förpackningsdirektivet , där denna kompromiss om att dela lika står , kan man se att detta inte fungerar .
förpackningar är fortfarande ett stort nedskräpningsproblem i europa och en belastning på miljön .
en del av socialisterna under ledning av bernd lange säger : &quot; ja , den här principen är bra , men vi skall inte införa den förrän år 2010 eller år 2012 enligt ändringsförslag 45 . &quot;
i den gemensamma ståndpunkten står det år 2006 .
enligt gruppen de gröna ger det bilindustrin mer än tillräckligt med tid att förbereda sig .
jag uppmanar därför mina kolleger att inte stödja kristdemokraternas ändringsförslag 38 och 45 av ett antal socialister .
om fordonstillverkarna själva måste stå för kostnaderna för återvinning av sina bilar , då kommer de att konstruera dem så att de blir lättare och billigare att återanvända .
då kommer problemet med plast , pvc , att försvinna från bilar och ersättas av bioplast framställd av växter .
när allt kommer omkring är det billigare , också för konsumenterna .
i tjugo års tid har en majoritet i parlamentet försökt att göra den europeiska miljöpolitiken grönare .
i dag hotar denna gröna position att gå förlorad under tryck från framför allt den tyska och franska bilindustrin .
därför , kolleger , rösta emot ändringsförslagen 38 och 45 .
vi i gruppen de gröna stöder i stora drag den gemensamma ståndpunkten .
herr talman ! avfallet från uttjänta bilar är ett av våra riktigt stora miljöproblem , både vad gäller avfallsmängd och utsläpp av miljöskadliga ämnen .
vi i gue / ngl-gruppen vill därför ha ett så heltäckande och konsekvent regelverk på området som bara är möjligt .
med detta direktiv har vi en möjlighet att ta ett stort steg framåt , men det förutsätter att rådets ståndpunkt inte trasas sönder och försvagas i parlamentets behandling .
flera av de ändringsförslag som har lagts fram skulle , om de antogs , försvaga direktivet mycket kraftigt .
det gäller framför allt ändringsförslag från ppe-gruppen , men tyvärr också några ändringsförslag från lange , som jag ser det .
det är inte svårt att ana att vissa länders bilindustri , t.ex. den tyska , har utfört ett ganska hårt lobbyarbete inför antagandet av detta direktiv .
för oss är det avgörande att följande principer skall gälla :
förorenaren skall betala .
det innebär att det är tillverkaren som skall ta det fulla ansvaret också ekonomiskt för återvinning av fordonen .
det måste finnas regler även för befintliga fordon .
vad gäller det kan vi inte godta att rådets ståndpunkt vad gäller datum för ikraftträdande skulle försvagas .
procentsatserna och kraven på återvinning vid vissa årtal får inte försämras . dessutom är det viktigt att begränsa användningen av farliga ämnen som bly .
vi kommer att rösta emot alla ändringsförslag som går i motsatt riktning i förhållande till detta .
om de ändringsförslag skulle antas som kraftigt försvagar direktivet , vore det mycket negativt , inte bara ur miljösynpunkt utan också för europaparlamentets trovärdighet i miljöfrågor .
det hänvisades tidigare i debatten till att man skall tänka på de miljoner människor som arbetar i bilindustrin i olika länder och de länder som har en stor bilindustri , t.ex. mitt eget hemland sverige .
jag har själv varit bilarbetare innan jag blev invald .
jag tror mig vara en av få i detta parlament som har stått vid ett löpande band och monterat bilar .
jag tycker att man skall ställa mycket hårda krav på bilindustrin .
det gynnar nämligen de moderna biltillverkarna som tänker miljövänligt och går snabbt framåt .
det är precis den typ av bilindustri som vi skall uppmuntra i europeiska unionen .
herr talman ! det gläder mig mycket att parlamentet nu prioriterar miljöskyddet , vilket medborgarna i europa med all säkerhet också gör .
det råder inget tvivel om , att övergivna bilar utgör ett allvarligt hot mot den visuella och fysiska miljön .
våra medborgare förväntar sig i detta hänseende att vi skall bevaka deras intressen .
varje år skrotas mellan 8 och 9 miljoner fordon inom europeiska unionen .
detta genererar i sig en stor mängd avfall .
biltillverkare , underleverantörer och tillverkare av utrustning måste anstränga sig för att begränsa användningen av farliga ämnen och måste därför i planeringsskedet se till att återanvänt material kan användas i tillverkningen av bilar .
vi vet att det i nederländerna finns auktoriserade behandlingscentraler som samlar upp uttjänta fordon , och denna metod bör spridas över hela europeiska unionen .
sett ur ett irländskt perspektiv vet jag att det irländska miljödepartementet redan har börjat samråda med företrädare för motorindustrin för att se till att lämpliga uppsamlingsplatser upprättas inom en snar framtid för att ta hand om uttjänta fordon på irland .
jag ser inget skäl till varför man inte skulle kunna organisera ett tillståndssystem för uppsamlingsplatser över hela europa , för att skrota de 8 till 9 miljoner fordon som man årligen gör sig av med inom europeiska unionen .
biltillverkare skall lämna information om hur stor del av de begagnade bilarna som kommer att kunna återanvändas , återvinnas och återställas under de kommande åren .
i enlighet med de nya bestämmelserna i amsterdamfördraget har samtliga 370 miljoner konsumenter inom europeiska unionen rätt till konsumentrelaterad information .
jag tror att eu : s konsumenter kommer att stödja de biltillverkare som tillämpar de miljövänligaste metoderna under det kommande året .
den sista frågan jag vill ta upp är att man i bestämmelserna och lagstiftningen måste ta hänsyn till den traditionella bilsektorns speciella ställning i hela den europeiska gemenskapen , på grund av den roll denna har i förhållande till den sociala sektorn samt mot bakgrund av miljömässiga och ekonomiska hänsynstaganden .
herr talman , ärade ledamöter ! direktivet om uttjänta fordon är verkligen en milstolpe på vägen mot en bättre miljö i detta vårt europa .
det verkar också som om man verkligen har ansträngt sig för att komma fram till en intelligent återanvändning av materialen , en minskning av det förorenande avfallet och ett främjande av tekniska innovationer .
vad detta beträffar är vi verkligen på rätt väg men , som några kolleger redan har betonat , är det reella problemet möjligheten att tillverkarnas ansvar blir ett solidariskt ansvar .
jag skulle vilja säga att man i italien har tagit betydande steg framåt på detta område . vi var kanske först i europa med att införa ett regelverk som uppmuntrar till att ta uttjänta fordon ur bruk , men vi har också i vårt land en ganska gammal bilpark och därmed allvarliga bekymmer för de marknadsproblem detta direktiv skulle kunna medföra .
jag tror att man måste analysera fenomenet på allvar .
i italien har man kommit till en inlämnings- och återvinningsgrad på omkring 80 procent , men det finns ett marknadsproblem som skulle kunna orsaka en smärre kris vad sysselsättningen beträffar . eftersom vi i italien har en industri som ofta tillgriper tillfälliga och permanenta friställningar kan detta medföra allvarliga svårigheter för löntagarna i olika delar av landet .
jag märker att parlamentet ibland är litet extremistiskt och intar ståndpunkter som antingen är ytterligt gröna eller raka motsatsen . därför tycker jag att man borde försöka förena de två kraven och finna en syntes .
resultatet är dessa intressanta ändringsförslag . här tror jag att man kan hitta en avvägd lösning på problemet , det vill säga att förena miljökraven med marknadens och sysselsättningens behov .
herr talman ! detta direktiv behandlar det förhållandevis lilla men växande problemet med övergivna bilar samt frågan om en mera strukturerad skrotning av uttjänta bilar .
i den utsträckningen kan det tänkas vara önskvärt , trots att det inte är något brådskande ärende .
huvudfrågorna är nu vem som betalar 262 euro per bil för de 9 miljoner bilar som skrotas varje år .
vem betalar för uppsamlingen , demonteringen , skrotningen och så vidare ?
och skall direktivet retroaktivt omfatta varje bil som någonsin tillverkats ?
kommissionens förslag , den allmänna ståndpunkten , är att tillverkarna skall betala allt .
detta skulle betyda miljarder pund eller euro för vart och ett av de större företagen i varje land inom europeiska unionen .
denna kostnad skulle ofrånkomligen föras över på priset och följaktligen på de nya bilarnas köpare .
eftersom europeiska biltillverkare har verkat här under många fler decennier än företag från japan , korea och andra länder , skulle det ligga till mycket större last för de äldre europeiska företagen och utgöra en konkurrensfördel för deras konkurrenter från andra länder .
jag uppskattar florenz , lange och andra som från partisplittringens båda sidor försökt uppnå en kompromiss baserad på delade kostnader .
jag rekommenderar också det ändringsförslag som jag undertecknat samt uppmanar mina kolleger från tyskland , italien , irland , spanien , sverige och storbritannien att eliminera denna åtgärds retroaktiva drag .
retroaktiv lag är dålig lag , den är ofta orättvis och ofta ogenomförbar .
de flesta demokratiska parlament i den fria världen förkastar den av princip såvida det inte föreligger ett överväldigande offentligt intresse , vilket det tydligen inte gör i det här fallet .
det är därför jag har manat till en omröstning med namnupprop om detta .
vi kan då se vem som är beredd att rösta för retroaktivitet med tvivelaktig legalitet , vilket skulle innebära en kostsam belastning för varje framtida bilköpare och ett förödande slag mot den europeiska bilindustrin .
herr talman , mina kära kolleger ! jag vill än en gång helt kort påminna om vilka ekonomiska frågor som står på spel med detta direktiv , och förnya mitt stöd till de ändringsförslag som min kollega bernd lange har ingivit .
fördelen med dessa ändringsförslag - jag vill insistera på detta - är att de sammanjämkar miljökrav och ekonomiska absoluta krav .
rådets gemensamma ståndpunkt innebär att biltillverkarna skall stå för hela eller en avsevärd del av kostnaderna för återtagande och återvinning av fordon .
men som lange så väl uttryckte det : för de europeiska tillverkarna är den lösningen fullkomligt orättvis .
eftersom jag kommer från ett land där det faktiskt finns biltillverkare , kan jag tala om att det är en omöjlighet att retroaktivt ålägga dem ett totalt finansiellt ansvar för alla de fordon som kommer från deras fabriker och som nu rullar på vägarna , vilket innebär ett ansvar för kostnader som ålagts 80 procent av den europeiska bilparken .
denna lösning är oacceptabel , eftersom tillverkarna inte har kunnat integrera miljökraven i sina tillverkningsprocesser och självkostnadspriser , de miljökrav som vi ålägger dem i dag .
den gemensamma ståndpunkten sätter de europeiska tillverkarna i ett ofördelaktigt läge gentemot de tillverkare som nyligen trätt in på den europeiska marknaden .
vi är självklart inte här för att försvara det ena eller andra nationella intresset eller den ena eller andra industrilobbyisten .
vi är däremot här för att bygga upp ett europa som kan konkurrera på världsmarknaden och för att försvara sysselsättningen inom de ekonomiska sektorer där vi faktiskt är konkurrenskraftiga .
av det skälet , kära kolleger , ber jag er att stödja de ändringsförslag som ingivits av bernd lange och som kommer att stödjas av europeiska socialdemokratiska partiets grupp .
faktum är att dessa ändringsförslag förlikar samtliga intressen - ekonomiska intressen och miljökrav - samtidigt som medlemsstaterna förblir fria att besluta om de närmare bestämmelserna för genomförandet av dessa krav , eftersom de system som nu gäller i medlemsstaterna - och det finns de som fungerar helt tillfredsställande - enligt förslagen skall få finnas kvar i fortsättningen .
herr talman , fru kommissionär ! det förslag till direktiv om uttjänta fordon som vi i dag ägnar oss åt syftar dels till att garantera ett starkt miljöskydd inom unionen , och dels till att säkra en fortsatt väl fungerande inre marknad för denna sektor .
jag vill bara kort säga att historiska bilar och veteranbilar givetvis skall undantas från tillämpningsområdet för detta direktiv .
vi är väl alla överens om att bilarna också utgör en del av vårt kulturarv .
en av stötestenarna avser artikel 12 , dvs. när direktivet skall börja tillämpas .
parlamentets föreslagna lösning , nämligen 18 månader efter det att direktivet trätt i kraft för nya bilar , är föga realistiskt .
den europeiska bilparken omfattar tiotals miljoner bilar som skall återtas utan att de har tillverkats för att återvinnas .
den gemensamma ståndpunkten var mer praktisk , eftersom den fastställde år 2006 för de bilar som redan är i trafik .
detta skulle dessutom ge företagen tid att uppbringa resurser för att hantera de tillkommande kostnaderna .
i likhet med min grupp kommer jag således att stödja den gemensamma ståndpunkten , som förefaller vara en balanserad kompromiss mellan företagens begränsningar och nödvändiga framsteg på miljöskyddsområdet .
herr talman , kära kolleger ! europaparlamentet står i dag inför ett viktigt beslut .
skall vi arbeta för ett framtidsorienterat miljö- och konsumentskydd eller skall parlamentet , vilket man kan befara enligt ändringsförslagen från florenz , lange och andra , göra sig till bödelsdräng åt den tyska bilindustrin ?
parlamentets trovärdighet som en av pionjärerna för miljöskydd står på spel .
det vore mer än genant om europaparlamentet skulle urvattna det som regeringarna i de 14 medlemsstaterna och europeiska kommissionen har beslutat vad gäller tillverkaransvaret och skyddet av miljön !
den avsikt florenz och lange har med ändringsförslagen är tydlig : direktivet skall förstöras !
genom det föreslagna delade ansvaret skall principen om att förorenaren skall betala urholkas och produktinnovationer undergrävas .
genom uppbyggnaden av talrika hinder vill de ingenting annat än att förhindra en effektiv ekologisk politik för avfallsströmmar , och via typgodkännanden vill de fördröja tillämpningen av direktiven med tolv år eller mer .
jag vädjar därför alldeles särskilt till de tyska ledamöterna : förhindra att det i dag uppstår en stor politisk skada !
den rödgröna förbundsregeringen har inte precis skördat några större lagrar i debatten om direktivet för uttjänta fordon .
låt inte detta fortsätta !
det ständiga gnället om konkurrensnackdelen är löjeväckande när det egentligen bara handlar om en konkurrensnackdel för den tyska bilindustrin .
var företrädare för folket , och låt er inte degraderas till företrädare för volkswagen !
rösta för miljö- och konsumentskyddet och för innovationer i bil- och återvinningsindustrin !
herr talman ! vi har diskuterat detta direktiv sedan 1997 .
nu är det dags att vi kommer fram till en överenskommelse .
eftersom jag mer eller mindre delar de åsikter som min kamrat sjöstedt och de grönas företrädare de roo framförde , tänker jag inte använda de två minuter jag har till mitt förfogande utan bara betona två frågor .
för det första , och det är kanske det viktiga i förslaget : tanken både angående återvinning och återanvändning om att man skall använda material som är mindre förorenande .
en annan viktig punkt är att avfall inte skall brännas eller sönderdelas , men inte bara när det gäller det som innehåller bly , kadmium och kvicksilver utan också det som innehåller pvc .
vi diskuterar denna fråga i ett annat forum i parlamentet .
den andra frågan gäller vem som skall stå för kostnaderna .
jag håller med de tidigare talarna när de säger att den som förorenar skall betala , och det har aldrig sagts bättre tidigare än i detta förslag .
tillverkarna skall betala , även om vi alla vet att kostnaderna i slutändan kanske läggs på konsumenterna , och de skall ta hand om kostnaderna före 2006 så som föreslås i vissa ändringsförslag .
vi instämmer mer med ändringsförslaget från första behandlingen .
det är också viktigt att fastställa en viss procent och det datum då fordonen skall bestå av återvinningsbart material .
jag tycker att man enligt förslaget förlitar sig på alltför långa tidsfrister .
slutligen , herr talman , anser jag att det är nödvändigt att gynna små och medelstora företag som , efter sträng kontroll och erhållande av vederbörliga tillstånd , kan skapa sysselsättning i detta så viktiga arbete , och på så sätt undvika storföretagens monopol .
herr talman , kära kolleger ! i dag måste europaparlamentet åta sig ett verkligt ansvar .
det handlar om vad vi skall göra med de miljoner fordon som vi överger varje år .
i vissa av våra stater har frivilliga miljöavtal redan tecknats för att våra diken , kanaler och fält inte längre skall fyllas av anskrämliga och farliga vrak , som en och annan skrämd höna har flytt .
jag kommer från ett land som är stolt över sin bilindustri och dess kommersiella framgångar , såväl i europa som i tredje land .
mitt lands internationella nimbus är en mätare på dess betydelse .
jag känner till den europeiska bilindustrins aktiva beteende ; den har satt igång ett omfattande forskningsprogram i syfte att upprätta ett nationellt informationssystem för nedmontering av gamla fordon .
jag är medveten om vilka svårigheter rådet har stött på för att finna en kompromiss .
därför måste vi i dag vara alkemister med förståelse och omsorg om vår miljö .
detta sekel kommer att bli avfallshanteringens sekel , i annat fall blir det inget sekel alls .
för min del bör man tillämpa principen att den som förorenar skall betala .
jag är säker på att bilindustrin , som visar en ständigt större respekt för miljön , har förväntat sig en sådan insikt .
den tar dessutom sitt ansvar .
men det åligger staterna att genomföra detta direktiv , och vi får akta oss för att göra det alltför detaljerat , eftersom de industriella traditionerna , nedmonterings- och skrotningsprocesserna ser olika ut beroende på om man är i italien eller finland .
jag motsätter mig det faktum att bilägarna skall göras ansvariga .
alla dessa kvinnor och män som rör på sig överallt i europa , de betalar sin bil , sin nationella skatt , sin katalysator , sin bränsleskatt - de betalar således redan ett mycket högt pris för denna fantastiska maskin och friheten att förflytta sig .
det skulle vara väl oförsiktigt - av mina kolleger i de stora grupperna med federalistisk böjelse - att vilja göra europaparlamentet så impopulärt genom att kunna tänka sig ett delat ansvar mellan ägaren och tillverkaren .
hur skall man dessutom kunna skapa en fond för att betala fordonsåtervinningen och förvaltningen av inomeuropeiska operationer ?
vem kommer att betala återvinningen av min bil som jag köpt i frankrike om jag låter registrera den i belgien ?
vilken nationell fond kommer att ta på sig ansvaret för mitt uttjänta fordon ?
vi får också akta oss för att oroa företagarvärlden med den rättsliga osäkerhet som har att göra med en oacceptabel retroaktivitet .
det är inte vår sak , här , att i dag dra igång en vedergällningsaktion med stöd av lagstiftning , vi bör i stället fortsätta på vår väg genom att förorda en hållbar utveckling .
herr talman ! europaparlamentet med utskottet för miljö , folkhälsa och konsumentfrågor i täten föresätter sig mestadels att kritiskt bedöma förslag från europeiska kommissionen eller rådet och förbättra dem från miljösynpunkt .
nu hotar en gedigen gemensam ståndpunkt från rådet att här i parlamentet bli sämre från miljösynpunkt .
varje år skrotar vi ett stort antal bilar med många farliga ämnen .
därför är förebyggande åtgärder med avseende på avfallsämnen viktiga .
vi bör också sträva efter så små mängder som möjligt av tungmetaller och andra farliga ämnen och material .
dessutom bör biltillverkarna ta hänsyn till att dessa bilar tillverkas på ett sådant sätt att det är enkelt att demontera och återanvända dem .
resterna av bilvraket kräver också en adekvat behandling .
jag stöder därför helhjärtat de procentsiffror för återanvändning och återvinning som föreslagits av rådet .
numera är det ekonomiskt möjligt att genomföra en fullständig demontering av bilvrak .
detta innebär att vi överger sönderdelning av bilvrak .
de uppställda målen är säkert genomförbara , och i nederländerna har återvinningen redan uppnått ett värde på 86 procent .
det bästa sättet att sörja för en god insamling är att den sista användaren kan lämna in bilen utan kostnad till en auktoriserad behandlingsanläggning .
kostnaderna för behandlingen kan sedan tas ut på priset för nya bilar .
de förslag som lagts fram av vissa parlamentsledamöter skadar detta system på ett allvarligt sätt .
det så kallade delade ansvaret är mycket opraktiskt och stimulerar inte till någon innovation .
om systemet med kostnadsfri inlämning tillämpas kommer det också att visa sig att kostnaderna för behandling kommer att sjunka avsevärt .
slutligen måste detta direktiv träda i kraft så snabbt som möjligt .
ett segdraget förlikningsförfarande innebär en onödig försening som går ut över miljön .
låt oss vara nöjda med den gemensamma ståndpunkt som nu föreligger ; då behöver vi inte göra någonting annat än att komplimentera och lyckönska rådet till det uppnådda resultatet .
herr talman ! jag vill ge kollega florenz ett stort erkännande .
han har under tryck , inte bara från sina kolleger utan också från bilindustrin , gjort ett gott arbete .
lägg därtill att florenz också var tvungen att göra detta med sin ekologiskt gröna inställning , var tvungen att mot den bakgrunden finna en kompromiss , och det var inte lätt .
allmänt sett är jag inte missnöjd med den gemensamma ståndpunkt som här ligger framför oss , och i vilket fall som helst inte med den filosofi som ligger bakom den gemensamma ståndpunkten .
det är två punkter som jag skulle vilja säga något om .
det gäller veteranbilarna och motorcyklarna , vilka mycket riktigt skall undantas från direktivet , och den andra punkten är hela den kontroversiella frågan om vem som egentligen bär ansvaret för återtagandet av bilarna .
jag vill inte tumma på texten i den gemensamma ståndpunkten .
producenten är ansvarig , måste vara ansvarig , och slutanvändaren måste utan kostnader kunna återlämna bilen .
jag tror att det finns för mycket ogrundad rädsla .
billobbyn har fört för många bakom ljuset .
jag vill därför än en gång säga till kollegerna att erfarenheterna visar att kostnaderna för denna behandling läggs på priserna .
det är inte så höga kostnader .
i den medlemsstat som jag kommer ifrån handlar det om 150 gulden per bil .
det innebär att man börjar på dag noll , och man kan då också behandla de gamla bilarna direkt .
då kan också en mycket stor industri direkt byggas upp som innebär att man ser till att de bilkyrkogårdar som tidigare var en vanlig syn i våra medlemsstater upphör att existera .
jag vill alltså inte tumma på den punkten i kompromissen .
jag tror att det är bra att vi så snabbt som möjligt sinsemellan godkänner den lagstiftning som nu ligger framför oss .
det är bra , eftersom det innebär att de nio miljoner bilar som varje år kommer ut på vägarna i europa också tas om hand på ett ordentligt sätt . det kommer oss allesammans till godo .
herr talman ! det föreliggande direktivet är en viktig åtgärd för att förebygga att vi får farligt avfall från uttjänta fordon , och det är viktigt för att främja återanvändning och återvinning av material från skrotade bilar .
jag menar därför att det är miljömässigt avgörande att förbudet mot att använda giftiga tungmetaller genomförs fullt ut , och att vi inte försvagar tillverkarnas ansvar .
gör vi detta tar vi bort incitamentet för tillverkarna att konstruera och tillverka bilar som ger mindre avfall .
det gemensamma systemet som efter mycket bekymmer antogs av rådet , som kommissionen stöder , och som också stöds av parlamentets utskott för miljö , uppfyller fullständigt de fastställda miljökraven och jag tycker därför att det är mycket egendomligt och oförståeligt att se ändringsförslag från ledamöter av utskottet för miljö som syftar till att väsentligt minska biltillverkarnas ansvar .
om dessa ändringsförslag antas , menar jag att parlamentets trovärdighet i miljöfrågor allvarligt måste ifrågasättas .
vi i parlamentet har hittills varit en positiv katalysator för miljöskydd och nu blir vi en negativ miljöfaktor i denna fråga i europa , om ändringsförslagen från florenz och lange antas .
om vi dessutom försvagar tillverkarnas ansvar i denna fråga , kommer det att få allvarliga konsekvenser för senare frågor på andra områden , t.ex. det kommande direktivet om elektronik- och datorskrot .
jag vill därför gärna uppmana parlamentets ledamöter att vi utan hänsyn till grupptillhörighet röstar emot alla de ändringsförslag till den gemensamma ståndpunkten som kommer att försvaga den miljömässiga standarden och som kommer att minska tillverkarnas ansvar .
på så sätt kan vi uppnå ett miljömässigt anständigt resultat .
herr talman ! detta förträffliga direktiv kommer att göra slut på dumpandet av gamla bilar , gynna återvinningen och framför allt uppmuntra tillverkarna att utforma bilar som lätt kan återvinnas .
men vem skall stå för kostnaderna ?
vilket system som än införs , kommer kostnaden slutligen att föras över på konsumenten .
det bästa sättet för oss att uppnå våra miljömål är att göra tillverkarna till vårt verktyg såväl för insamlingen av pengarna som för skrotningen och återvinningen av bilarna .
tillverkarna har lurat florenz och lange att lägga fram ändringsförslag här som allvarligt försvagar dessa förslag .
låt er inte luras av biltillverkarna !
om ni vill dra full nytta av detta direktiv , använd er röst till att förkasta dessa ändringsförslag .
herr talman , fru kommissionär , kära kolleger ! i motsats till vad vi skulle kunna tro är denna debatt inte av teknisk art .
den har blivit högst politisk .
i går hedrade vi vår institution med en politisk debatt - vi skulle vanhedra oss själva om 314 ledamöter i dag gav efter för vissa biltillverkares lobbygrupper .
genom att begära att konsumenterna skall stå för hälften av kostnaderna för återtagande av uttjänta fordon , vilket ändringsförslag 38 föreskriver , samtidigt som den gemensamma ståndpunkten kräver att tillverkaren skall ansvara för hela återtagandet , skulle europaparlamentet för första gången inte framträda som en garant för försvaret av de europeiska konsumenterna och medborgarna , utan i stället bli något av en resonanslåda för lobbygrupperna .
det skulle vara ett prejudikat som öppnade dörren för alla slags påtryckningar inom många andra områden .
det skulle också vara första gången som europaparlamentet försvagade rådets ståndpunkt , när vi i allmänhet kritiserar rådets ståndpunkter för att inte räcka till .
ett system för gratis återtagande av gamla fordon och ett utökat antal fordon som skall återvinnas är exempel på åtgärder som kommer att få såväl återvinningsverksamheten som den därmed förknippade sysselsättningen att växa .
med tanke på konsumenterna , miljön och de nya arbetstillfällen som kan skapas inom återvinningssektorn , får vi absolut inte ändra rådets gemensamma ståndpunkt , som i sin nuvarande version är helt godtagbar .
herr talman ! liksom så många andra här i dag tror jag att detta är en bra åtgärd .
det är en nyttig åtgärd och nödvändig för oss alla .
de flesta tekniska frågorna är lösta .
det återstår att slutgiltigt godkänna vissa detaljer , men de flesta tekniska frågorna är lösta .
vi har kommit fram till den sista frågan .
under debatten vid den första behandlingen var det endast utskottet för ekonomi och valutafrågor som ställde den här frågan och det var bara jag själv i egenskap av den som författat utskottets yttrande som ställde den frågan i parlamentet .
den är mycket enkel : vem betalar ?
kommissionens allmänna ståndpunkt innebär en rimlig kompromiss på så sätt att tillverkarna skall betala en betydande del av kostnaden , inte hela kostnaden som bowis nämnde av misstag .
i själva verket så litet som 20 procent eller en femtedel av kostnaderna , enligt juristerna .
detta är inte orimligt .
om man ser på konsumenten i storbritannien som köper en rover , som lange pekat på , eller vilket annat bilmärke i storbritannien som helst för den delen och som i åratal har betalat överpriser för dessa bilar , långt över jämförbara priser i andra delar av europa , varför skall de betala ?
de har redan betalat .
varför skulle de här människorna , som skattebetalare eller som framtida bilköpare , åter betala för skrotning av ett fordon som tillverkaren har gjort vinst på ?
jag kan inte acceptera det .
enligt vissa ändringsförslag här i dag föreslås det att detta bör vara fallet .
jag kan inte acceptera det och jag kommer inte att rösta för det .
ansvaret för dessa bilar ligger hos tillverkaren .
det är tillverkaren som måste sörja för infrastrukturen och stå för en rimlig del av skrotningskostnaderna .
den gemensamma ståndpunkten utesluter inte möjligheten att staten skulle kunna ge bidrag .
den gemensamma ståndpunkten är en rimlig kompromiss .
en del av dagens ändringsförslag är fullständigt orimliga då de helt och hållet fråntar biltillverkaren ansvaret för att betala en liten del , om ens någon , av skrotningskostnaden för bilar i användning .
jag kan inte acceptera detta och på skattebetalarnas och de europeiska konsumenternas vägnar röstar jag emot dessa ändringsförslag .
herr talman , mina ärade damer och herrar ! det råder enighet om att vi måste börja tänka på hur vi i europa skall handskas ordentligt med gamla bilar , men rådet har i detta fall inte gett något exempel på en meningsfull europeisk miljöpolitik .
det var blamerande hur det tyska ordförandeskapet behandlade frågan .
först stämde trittin , miljöministern , inte av det hela i tillräcklig utsträckning med sina kolleger i kabinettet , därpå kom förbundskansler schröder likt en elefant i en porslinsbutik och blandade sig utan sakkunskap i förfarandet .
men inte heller beslutet från det finländska ordförandeskapet i juni var det bästa man kunde uppnå . det finns ett par svagheter .
den största svagheten är som jag ser det att man inte har tagit tillräckligt stor hänsyn till de medelstora företagens situation , men bilindustrin består inte endast av storföretag .
just på underleverantörsområdet spelar medelstora företag en mycket stor roll , och vi måste ta hänsyn även till de anställdas intressen i dessa små och medelstora företag .
därmed är det långt mer än två miljoner människor som har sitt arbete på detta område .
många ändringsförslag från utskottet för miljö , folkhälsa och konsumentfrågor gagnar just de medelstora företagen , liksom också de föreliggande ändringsförslagen från vår grupp till artikel 5 gällande kostnaderna .
inte heller från miljöpolitisk synpunkt är den gemensamma ståndpunkten någon lysande prestation .
det saknas blick för de stora sammanhangen , och när kollegan från de gröna säger att det skulle bli första gången som europaparlamentet försvagade den gemensamma ståndpunkten så är det ingenting man kan påstå , för ur ett miljöpolitiskt perspektiv är det ju föga meningsfullt om vi genom stela , höga återvinningsmål hindrar moderna , energisnåla fordon såsom 3-liters-bilen , där det ju används mycket plast !
därför måste man stödja ett ändringsförslag som innebär att man åtminstone tolererar undantag om vi har särskilt sparsamma bilar .
industrins invändningar är säkerligen inte ologiska på detta område .
plast- och bilindustrins argumentationskraft skulle emellertid tillta även om man inte bara i detta sammanhang skulle engagera sig för en reducering av koldioxid i europa .
herr talman ! i dag befinner vi oss verkligen i en ovanlig situation : de som vill försvara miljövärdena ställer sig bakom rådets gemensamma ståndpunkt .
till skillnad från föregående talare kan jag konstatera att jag verkligen är stolt över att man under det finländska ordförandeskapet kom fram till en gemensam ståndpunkt som försvarar miljövärdena .
om vi frångår den gemensamma ståndpunkten och strävar efter att dela kostnaderna för återvinning skapar vi kryphål : vi får inte något vettigt , klart system där ansvarsförhållandena är i sin ordning .
därför är det enligt min mening tillverkaren som skall bära huvudansvaret .
det är bara så vi kan lösa problemet på ett tillräckligt bra sätt och även ta hänsyn till att tillverkarna uppmuntras att tillverka sådana fordon som i framtiden kan återvinnas till så låga kostnader som möjligt .
herr talman ! det finns två principiella frågor i rådets förslag till direktiv .
den ena rör producentens oinskränkta ansvar att återta uttjänta fordon .
det riskerar att det skapas en monopolsituation inom demonteringsverksamheten .
särskilt gäller detta i områden inom eu där avstånden är stora , och där många småföretag är engagerade i demontering .
jag menar att eg : s direktiv inte får , oavsett vad ärendet gäller , missgynna de små företagen inom unionen .
producenternas oinskränkta ansvar riskerar även att marknaden för begagnade bildelar försvinner . en producent har ett större ansvar att sälja nya delar .
denna handel är viktig , särskilt för dem som samlar på och renoverar äldre fordon .
denna princip är även tveksam utifrån marknadsekonomiska principer .
företag skall kunna förändras , säljas och avvecklas .
de skall kunna etablera sig på nya marknader , men även lämna gamla marknader .
att binda producenter med ett ansvar som kan sträcka sig mycket långt bakåt i tiden stämmer illa med en flexibel och utvecklingsfrämjande marknadsekonomi .
den andra principen i rådets gemensamma ståndpunkt är inslaget av retroaktivitet i direktivförslaget .
det strider mot vedertagna ekonomiska och juridiska principer , att retroaktivt ålägga en producent ekonomiskt ansvar för sin vara .
det ändrar även ägaransvaret retroaktivt .
en konsument kan under åren ha ändrat produkten i flera avseenden .
alla länder inom eu har i dag lagar som reglerar skrotning av bilar .
de kan vara bättre och de kan vara sämre länderna emellan .
i avvaktan på att detta eg-direktiv får genomslag bör emellertid eu-länderna , var för sig , ansvara för skrotning av fordon på bästa sätt , så att retroaktiviteten i eu-lagstiftningen inte tillämpas .
detta strider inte mot en finansieringsmodell med fonduppbyggnad .
herr talman ! att den åtgärd vi diskuterar är viktig för miljön och industrin är uppenbart och någonting vi alla kan enas om .
den gemensamma ståndpunkten är en godtagbar men mycket känslig och vansklig kompromiss , så mycket mer eftersom den medför ganska begränsade förbättringar om man inte skall äventyra hela direktivet .
jag hävdar alltså att parlamentet inte kan utöva tvång och att det vore paradoxalt om det skulle göra det om en linje som innebär en minskning av åtgärdens miljökonsekvenser .
jag påminner om att biltillverkarna har medgett att de kan leva med direktivet . kostnaderna är inte astronomiska : att återvinna en bil kostar mindre än 1 procent av nybilspriset .
dessutom träder tillverkarnas ekonomiska ansvar inte i kraft förrän år 2006 , när en stor del av dagens fordonspark inte längre finns på marknaden .
för de återstående fordonen kan man också införa en slags ansvarsfördelning , såsom föreslås i langes ändringsförslag 44 och 45 , de enda jag tycker är förenliga med balansen i den gemensamma ståndpunkten och med de aktuella erfarenheterna i somliga länder , och som därför är värda att stödja .
herr talman ! detta är ett ytterst dåligt direktiv .
för det första , som min kollega bowis har påpekat , är det retroaktivt och därför principiellt felaktigt .
för det andra , det lägger enorma kostnader på den europeiska fordonsindustrin , vilket skulle skada konkurrenskraften och sysselsättningen .
i det här parlamentet diskuterar vi ständigt behovet av att främja sysselsättning och arbetstillfällen i europa och ändå vidtar vi ständigt åtgärder som kommer att ha ett negativt inflytande på sysselsättningen .
jag vill påstå att direktivet är dåligt även i ett annat avseende , vilket inte har granskats tillräckligt grundligt i denna debatt .
det är som mycket annat i europeisk lagstiftning .
det är alldeles för normativt .
det cementerar en specifik återvinningsmodell .
det löpande bandet uppfanns för cirka hundra år sedan , jag tror det var av henry ford , och det som vi håller på att göra här övertygar mig om att vi försöker skapa något slags omvänt löpande band i artonhundratalsstil - för att demontera fordon , för att ta isär delarna och försöka återvinna dem .
en sak som vi borde tänka på är att marknaden för återvunna stötfångare i plast är mycket osäker .
plastindustrin vill för det mesta inte ta tillbaka dessa delar och kan av ekonomiska skäl inte heller göra detta .
det finns redan en mycket framgångsrik industri som skrotar bilar , återvinner metaller och återvinner energi genom förbränning av icke-metalldelar .
detta är ett ur miljösynpunkt mycket rimligt tillvägagångssätt .
miljömässigt sett är det lika bra att bränna gammal plast som att bränna ny olja för energiåtervinning .
denna bilskrotningsmetod medför inga kostnader och skulle sålunda eliminera hela frågan om vem som betalar , eftersom den &quot; döda &quot; bilen i själva verket har ett lågt värde då den kommer in i återanvändnings- och återvinningsprocessen .
jag motsätter mig detta direktiv eftersom det är för normativt , det tar ingen hänsyn till vad som för tillfället i själva verket pågår på bilåtervinningsmarknaden , och det cementerar metoder som inte nödvändigtvis är de bästa ur miljösynpunkt och säkerligen är mycket skadliga ekonomiskt sett .
herr talman , kolleger ! den gemensamma ståndpunkten är bra , men det är parlamentets uppgift att ytterligare förbättra den gemensamma ståndpunkten om uttjänta fordon .
den socialdemokratiska gruppen har under de senaste dagarna kommit med några viktiga förslag till förbättring .
jag skulle framför allt vilja göra er uppmärksamma på ändringsförslag 45 . där väljer vi att lägga kostnaderna för demontering och återvinning hos producenterna , i alla fall för nya bilar .
i samband med konstruktion och produktion kommer man därigenom att ta hänsyn till återvinning .
för de bilar som nu är i trafik är det rimligt att dela kostnaderna , till exempel genom att inrätta en fond som i nederländerna .
i den gemensamma ståndpunkten står det att producenterna inte bara skall stå för kostnaderna , utan att de också måste ta tillbaka de uttjänta bilarna .
det är enligt min uppfattning ett mycket stort problem .
jag pläderar för att inte låta just biltillverkarna organisera skrotning och återvinning , för det skulle leda till att tillverkarna får ett för stort grepp om marknaden för begagnade delar .
de kan då själva bestämma priserna .
var och en som någon gång har kört en gammal bil vet att detta är till nackdel för konsumenten och för den som gillar att meka .
den europeiska konsumentorganisationen , som bett oss att stödja den gemensamma ståndpunkten på den punkten , lämnar enligt min mening konsumenten i sticket .
ett andra argument för att hålla bilskrotningen borta från tillverkarnas händer är transportkostnaderna .
om alla biltillverkare kommer att inrätta sina egna skrotningsföretag kommer det att göra det nödvändigt att bogsera bilvrak över långa avstånd .
det är både miljöovänligt och dyrt . inte heller detta har konsumenten någon nytta av .
därför skulle jag gärna se att ni stöder ändringsförslag 45 .
herr talman ! det förslag som vi diskuterar innehåller ett mycket stort antal positiva punkter , företrädesvis inriktade på att förebygga avfall , återanvändning , återvinning och recirkulation av delar , återvinning av material och så vidare .
jag tror att vi har lämnat ifrån oss ett bra förslag .
diskussionen handlar företrädesvis om ifall konstruktören , den slutliga försäljaren eller någon annan måste ta tillbaka bilvraket gratis eller inte .
jag skulle bara vilja ta mitt eget land som exempel för att förklara hur det fungerar där utan några problem .
vi har nått en överenskommelse med alla dem som berörs av denna fråga , det vill säga bilkonstruktörerna , de som handlar med begagnade bilar , bilindustrins samarbetsorganisation , behandlingsanläggningarna för metall , sönderdelningsanläggningarna och staten .
det finns ett miljöpolicyavtal som undertecknats på frivillig väg .
bilindustrin , och belgien är ett land med en mycket stor bilproduktion , har inte ställt till med något som helst problem i samband med detta .
våra medborgare kan lämna in sin bil gratis till den slutliga försäljaren .
tvärt emot vad som sägs här , om att detta skulle vara till nackdel för sysselsättningen , har vi kunnat konstatera hur en rad småföretag helhjärtat tagit sig an återvinningen av materialet , och att de gör det på ett mycket bra sätt .
vissa företag har blivit spetsföretag eftersom de lyckats återvinna vissa material , till och med material som ännu inte är upptagna i direktivet .
det innebär således att vi här utvecklar en ny sektor , ny sysselsättning och gör miljön en stor tjänst .
jag är för gratis inlämning .
det har lyckats hos oss .
varför skulle det inte kunna lyckas någon annanstans ?
herr talman , ärade parlamentsledamöter ! tack för en intressant debatt med många viktiga argument som har framförts .
vill ni vara snälla att stå ut med mig under att par minuter .
tillåt mig att kort redogöra för några av de utgångspunkter och principer som ligger bakom detta direktiv .
låt mig också börja med att kommentera och svara på ett par av de viktigaste argumenten i denna debatt .
för det första tror jag att vi skall upprepa några grundläggande fakta som redan florenz och andra har nämnt .
det vi diskuterar här är det faktum att närmare tio miljoner bilar skrotas varje år i europeiska unionen , att det utgör ungefär lika många miljoner ton avfall .
det vill säga närmare tio miljoner ton avfall skapas av dessa bilar , och ungefär 7 procent av dessa lämnas i naturen .
de utgör dessutom miljöfarliga ämnen av värsta slag .
ungefär 10 procent av produktionen av bly återfinns i bilar , men också kadmium , krom , kvicksilver och andra mycket farliga ämnen .
detta känner ni redan till , men jag vill ändå upprepa det också för dem som lyssnar .
detta är en av de snabbast växande avfallsströmmarna som vi har i europa .
vi vet att avfallet finns där , vi vet hur vi skall handskas med det , och det finns ingen ursäkt för att undvika att handla .
det finns tre syften med detta direktiv : för det första vill vi få bort användningen av giftiga tungmetaller från tillverkningen av nya bilar .
vi vill för det andra slå fast tillverkaransvaret .
vi kan inte längre ta hand om saker i slutet av en produkts livscykel , utan vi skall undvika att skapa så mycket av avfall .
vi skall se till att återvinna så mycket som möjligt av en produkts olika innehåll .
för det tredje vill vi nå återvinningsmål som är preciserade i detta direktiv .
det är de tre viktigaste syftena med direktivet .
det beror ju på att det är ett slöseri med resurser att vi inte ser till att materialet som finns i bilar återvinns .
det är framför allt producentens resurser som vi slösar med om vi inte tar itu med en bils livscykel .
två viktiga frågor har kommit upp här - ja , det finns fler , men jag vill nämna två av de viktigaste .
för det första : vem skall betala ?
den andra frågan är : försämrar vi europeisk bilindustris konkurrenskraft med detta förslag ?
den första frågan gäller alltså vem som skall betala .
i direktivet framgår det att kostnaden skall bäras huvudsakligen av producenten i enlighet med de principer som vi har i eu : s fördrag om producentansvar samt att förorenaren skall betala .
det är dock klart att denna kostnad kommer att bäras gemensamt av producenter och konsumenter .
vi har räknat ut att kostnaden för att återvinna bilar inte utgör mer än en procent av priset för en ny bil .
tror vi då att kostnaden försvinner , om vi inte skulle anta detta direktiv ?
nej , det är klart att vi alla kommer att få bära kostnaden för att miljön förstörs , men det blir mycket dyrare .
dessutom kommer kostnaden längre fram .
kostnaden försvinner alltså inte , men nu tydliggör vi vems ansvaret är och hur kostnaden skall fördelas .
talar vi då om en bilindustri i kris ?
är det en vinstsvag industri som vi diskuterar och som vi verkligen måste hjälpa genom att inte lägga på fler pålagor ?
är det så att bilindustrin absolut inte har råd ?
är det så att motiven i själva verket är att försämra europeisk bilindustris konkurrenskraft ?
det är alldeles tvärtom !
tror ni att konsumenternas krav på miljövänliga bilar och bränslesnålare bilar kommer att minska i framtiden ?
vad tror ni att barn och barnbarn kommer att ställa för krav på bilar , eller att lagstiftarna i framtiden kommer att ställa för krav på bilar ?
naturligtvis att de skall vara miljövänliga , att de skall kunna återvinnas , att de skall vara bränslesnåla , att de inte skall förorena vår miljö !
det är ju bara på detta sätt som vi kan skapa en framtid för bilindustrin .
vi måste skapa drivkrafter som är sunda , som ser till att vi tar hand om avfallet , att vi återvinner materialet , att vi kan konkurrera med miljövänliga och bränslesnåla bilar .
det faktum att vi har en europeisk bilindustri som redan är långt framme kompenserar mer än väl att det faktiskt finns fler bilar som de måste ta ansvar för , som rullar i europa .
detta är ingen oöverstiglig kostnad eller oöverstiglig uppgift .
om vi skapar sådana drivkrafter kommer - det är jag helt säker på - marknadskrafterna och de kommersiella intressena i bilindustrin att se till att det växer fram system för att ta hand om både det ena och det andra .
det kommer att bli allt från försäkringar till bra och vettiga skrotningssystem och återvinningssystem .
det kommer industrin själv att se till att det uppstår i europa .
detta är ingen oöverstiglig kostnad för europeisk bilindustrin .
det kommer i stället att hjälpa industrin att vara i fronten när det gäller att producera miljövänliga och bränslesnålare bilar så småningom .
detta måste vi göra för miljöns skull .
kostnaderna försvinner inte , avfallet försvinner inte .
annars måste vi alla som skattebetalare eller samhällsmedborgare betala notan ; dessutom blir det dyrare om vi gör det längre fram , ju längre vi väntar .
detta skulle jag vilja säga inledningsvis .
jag vill också kommentera frågan om det är retroaktiv lagstiftning .
om vi räknar med att en bil i genomsnitt lever elva år , menar parlamentarikerna , eller menar någon , att vi skulle vänta elva år framåt i tiden innan vi tar itu med detta problem ?
menar ni att vi när vi lagstiftar om kemikalier skulle säga att vi inte låtsas om de kemikalier som redan finns på marknaden , och att vi bara lagstiftar för det som skall tillverkas längre fram i tiden ?
det är klart att vi måste se på det problem som just nu finns där och den utmaning som den existerande bilparken utgör .
det är fortfarande inget oöverstigligt problem .
vi kan ta hand om det .
vi har redan en infrastruktur .
vi har det som vi behöver för att ta hand om uttjänta bilar .
jag hoppas naturligtvis att resultatet av omröstningen skall bli bra i dag .
jag vill också , om jag inte redan har gjort det , tacka karl-heinz florenz för det hårda arbete som han har lagt ned i miljöutskottet på detta förslag .
det är faktiskt i många avseenden banbrytande vad gäller återanvändning och producentansvar .
jag tror att det kommer att få mycket positiva och märkbara effekter på miljön .
vi kan inte fortsätta att blunda för det .
vi har som sagt både kunskaperna och tillgångar för att klara av detta .
efter den första behandlingen i europaparlamentet 1999 hamnade kommissionens förslag i en besvärlig politisk situation i rådet .
vi fick emellertid en väl avvägd gemensam ståndpunkt i juli under det finländska ordförandeskapet .
nu måste vi se till att denna lagstiftningsprocess avslutas på ett framgångsrikt sätt .
det har lagts fram sammanlagt 48 ändringsförslag .
kommissionen kan anta 10 ändringsförslag helt och hållet .
tre ändringsförslag kan godtas delvis , och ett kan godtas i princip .
vissa ändringsförslag rör förbättringar av kommissionens förslag som vi godtog redan vid den första behandlingen , eller återinför i direktivet sådana delar av det ursprungliga förslaget som rådet har tagit bort .
detta gäller ändringsförslag 5 , utom första delen , 8 , 9 , första delen , 10 , 12 , tredje delen , 15 , 16 , 20 , 22 , 24 och 25 .
dessa ändringsförslag kan alla godtas .
ändringsförslag 6 och 21 är nya ; kommissionen kan godta dem .
kommissionen kan också godta ändringsförslag 26 med vissa redaktionella ändringar .
jag vill betona att ett antal av de övriga ändringsförslagen som rör förslagets grundläggande komponenter innebär en avsevärd urvattning av den miljöskyddsnivå som är syftet med den gemensamma ståndpunkten .
de kan därför inte godtas .
parlamentet har av tradition starkt bidragit till att stärka miljölagstiftningen i europa .
det skulle förvåna mig och göra mig nedstämd om så inte blev fallet i dag .
jag är mycket bekymrad över vissa ändringsförslag från parlamentet som ifrågasätter det här förslagets absoluta grundpelare .
det rör t.ex. utfasning av tungmetaller , tillverkaransvaret och återvinningskravet .
jag vill bemöta dessa ändringsförslag gruppvis .
ändringsförslagen 4 , 11 , 12 , 13 , 28 , 30 , 32 , 37 , 42 och 48 gäller utfasningen av tungmetaller .
ändringsförslag 12 innebär att bestämmelsens ikraftträdande försenas med minst 10 år .
ändringsförslagen 13 , 28 , 32 , 37 , 42 och 48 innebär att onödiga villkor och undantag införs .
det skulle innebära att processen med att ersätta de skadliga ämnena kommer att gå långsammare .
ändringsförslagen 4 , 11 och 30 innebär att tungmetaller måste avskiljas från avfallet före återvinning .
kommissionen anser att den utfasning som föreslås i den gemensamma ståndpunkten är lättare att tillämpa ur teknisk synvinkel .
ändringsförslagen 17 , 18 , 27 , 34 , 36 , 38 , 44 och 45 gäller tillverkaransvaret .
den kompromiss som rådet har kommit fram till är rättvis men skör .
kommissionen anser inte att ändringsförslagen skulle förbättra balansen utan att samtidigt skapa spänningar .
jag beklagar den förvirring som uppstod nyligen genom att interna dokument från kommissionen användes på fel sätt , vilket skapade ovisshet om kommissionens inställning i frågan .
jag vill betona att kommissionen redan 1997 föreslog en särskild klausul om tillverkaransvar , och att kommissionen helt stöder den gemensamma ståndpunkten .
det lägger inte oproportionerliga kostnader på tillverkarna , långt därifrån .
ändringsförslagen 39 , 40 , 46 och 47 gäller kvantifierade mål .
den höga skyddsnivå som den gemensamma ståndpunkten syftar till skulle urholkas mycket om återvinningsmålet för 2006 tas bort .
dessa ändringsförslag skulle också göra målen besvärliga att handskas med och svåra att övervaka .
låt mig dessutom kommentera - lyssna noga på vad jag säger nu , eftersom jag har hört detta upprepas i debatten - frågan om veteran- och hobbybilar som nämns i ändringsförslagen 3 , 7 , 9 , andra delen , och 35 .
sådana fordon omfattas inte av definitionen om avfall och omfattas därför inte av direktivet .
så vad som än har påståtts här omfattas inte veteranbilar och motorcyklar av direktivet .
vi anser inte att ändringsförslagen 2 och 14 tillför direktivet något .
ändringsförslag 23 innebär att kommissionen måste anta kvalitetsnormer för återanvändbara komponenter .
detta omfattas inte av direktivet .
det skulle därför krävas ett ad hoc-direktiv från europaparlamentet och rådet .
ändringsförslagen 29 , 31 och 41 urvattnar demonteringskraven .
särskilt ändringsförslagen 31 och 41 riskerar att urholka möjligheterna att återvinna plast , däck och glas .
kommissionen kan slutligen inte godta ändringsförslagen 1 och 33 av skäl som har med den rättsliga klarheten att göra samt ändringsförslag 19 som kommissionen anser vara onödigt på detta stadium .
ändringsförslag 43 hör vidare inte hemma i direktivets tillämpningsområde .
omröstningen kommer härefter att äga rum .
( en ) fru talman ! som ni vet är orsaken till att vi röstar om det här betänkandet i dag och inte i förra veckan de talrika översättningsfelen , särskilt i den franska versionen .
ni har fått en klagoskrivelse av mig angående antalet felaktigheter i detta betänkande samt i andra betänkanden som jag har haft att göra med på sista tiden .
ett fel som ännu inte har rättats till finns i ändringsförslag 4 .
i den engelska versionen avser vi farmakologiska och vetenskapliga organisationer .
i den franska versionen står det &quot; entreprises pharmaceutiques et organisations scientifiques &quot; .
kan ni vänligen se till att de fransktalande parlamentsledamöterna får veta att ordet entreprises inte är korrekt .
det skall inte finnas med i ändringsförslaget .
och jag ber er igen , fru talman , att se över standarden på de översättningar vi för närvarande får ta emot .
fru mcnally ! generellt sett är jag själv också bekymrad över att översättningarna ställer till med allt fler problem .
jag skall höra med enheterna om hur vi skall kunna lösa detta .
betänkande ( a5-0011 / 2000 ) av langen för europaparlamentets delegation till förlikningskommittén om förlikningskommitténs gemensamma utkast till europaparlamentets och rådets beslut om ett flerårigt program för främjande av förnybara energikällor inom gemenskapen ( 1998-2002 ) - altener ( c5-0333 / 1999 - 1997 / 0370 ( cod ) )
betänkande ( a5-0010 / 2000 ) av ahern för europaparlamentets delegation till förlikningskommittén om förlikningskommitténs gemensamma utkast till europaparlamentets och rådets beslut om antagande av ett flerårigt program för att främja en effektiv energianvändning ( 1998-2002 ) - save ( c5-0334 / 1999 - 1997 / 0371 ( cod ) )
betänkande ( a5-0009 / 2000 ) av graca moura för europaparlamentets delegation till förlikningskommittén om förlikningskommitténs gemensamma utkast till europaparlamentets och rådets beslut om att inrätta ett enhetligt instrument för finansiering och programplanering för kulturellt samarbete ( kultur 2000-programmet ) ( c5-0327 / 1999 - 1998 / 0169 ( cod ) )
andrabehandlingsrekommendation ( a5-0006 / 2000 ) för utskottet för miljö , folkhälsa och konsumentfrågor om rådets gemensamma ståndpunkt ( 8095 / 1 / 1999 - c5-0180 / 1999 - 1997 / 0194 ( cod ) ) inför antagandet av europaparlamentets och rådets direktiv om uttjänta fordon ( föredragande : florenz )
betänkande ( a5-0007 / 2000 ) av berger för utskottet för rättsliga frågor och den inre marknaden om förslaget till europaparlamentets och rådets direktiv om utstationering av arbetstagare från tredje land i samband med tillhandahållande av tjänster över gränserna ( kom ( 1999 ) 0003 - c5-0095 / 1999 - 1999 / 0012 ( cod ) )
betänkande ( a5-0012 / 2000 ) av berger för utskottet för rättsliga frågor och den inre marknaden om förslaget till rådets direktiv om en utvidgning av friheten att tillhandahålla tjänster över gränserna till att även omfatta tredjelandsmedborgare som har etablerat sig inom gemenskapen ( kom ( 1999 ) 0003 - c5-0050 / 2000 - 1999 / 0013 ( cns ) )
betänkande ( a5-0003 / 2000 ) av marinho för utskottet för rättsliga frågor och den inre marknaden om
i. förslaget till rådets beslut om ändring av beslut 88 / 591 / eksg , eeg , euratom om upprättandet av europeiska gemenskapernas förstainstansrätt ( 5713 / 1999 - c5-0020 / 1999 - 1999 / 0803 ( cns ) )
ii. förslaget till rådets beslut om ändring av beslut 88 / 591 / eksg , eeg , euratom om upprättandet av europeiska gemenskapernas förstainstansrätt ( 9614 / 1999 - c5-0167 / 1999 - 1999 / 0805 ( cns ) )
( genom på varandra följande omröstningar antog parlamentet de två lagstiftningsresolutionerna . )
betänkande ( a5-0022 / 2000 ) av brok för utskottet för utrikesfrågor , mänskliga rättigheter , gemensam säkerhet och försvarspolitik om förslaget till rådets beslut om exceptionellt finansiellt stöd till kosovo ( kom ( 99 ) 0598 - c5-0045 / 2000 - 1999 / 0240 ( cns ) )
fru talman ! jag skulle bara vilja påpeka att enligt förfarandet medges inte varken att man framlägger eller följaktligen röstar om ändringsförslag i utskottet .
jag vet inte om detta är enligt reglerna och därför uppmanar jag er att kontrollera om det förfarande som följdes innan denna åtgärd kom till kammaren var korrekt .
jag noterar det ni just sade , herr speroni .
betänkande ( a5-0018 / 2000 ) av dimitrakopoulos och leinen för utskottet för konstitutionella frågor om sammankallandet av regeringskonferensen ( 14094 / 1999 - c5-0341 / 1999 - 1999 / 0825 ( cns ) )
gemensamt resolutionsförslag om förhandlingarna om regeringsbildningen i österrike .
fru talman ! även på detta område har vi som vanligt ett antal översättningsproblem .
som utgångspunkt gäller den engelska versionen .
för att ge er ett exempel har det fallit bort något i såväl den nederländska som i den tyska versionen vid punkt 4 liksom vid punkt 5 , och jag citerar de fyra orden på engelska : &quot; in so far as &quot; .
jag skulle därför vilja be er att använda den engelska versionen som utgångspunkt .
tack , herr van velzen .
jag säger samma sak till er som jag sade till mcnally för en stund sedan .
jag är mycket bekymrad över de översättningsproblem som blir allt vanligare , och jag kan försäkra er att vi kommer att se på detta mycket , mycket allvarligt .
under alla omständigheter är det givetvis originalversionen som är den gällande .
. ( fr ) jag gläder mig åt detta utmärkta betänkande om meddelandet &quot; kvinnor och vetenskap &quot; !
i detta dokument föreslår kommissionen att vi skall stimulera debatten i syfte att främja kvinnors ökat deltagande i den europeiska forskningen .
det är ett mål som förtjänar allt vårt stöd .
utgifterna för forskning och teknik utgör en ansenlig del av europeiska unionens budget , efter jordbruket och strukturfonderna .
de olika ramprogrammen har inte endast möjliggjort vetenskapliga arbeten av hög kvalitet , utan också ett nydanande samarbete mellan forskare från olika medlemsstater .
samtidigt finns det få kvinnor inom de vetenskapliga disciplinerna , trots att de uppnår mycket goda resultat under sina studier .
kvinnornas underrepresentation får inte fortgå .
därför välkomnar jag med nöje europeiska kommissionens förslag .
syftet med detta dokument är en koncentration på åtgärder att vidta på gemenskapsnivå , och mera särskilt via det femte ramprogrammet för forskning och teknisk utveckling , något jag självklart stöder .
under de kommande åren gäller det att öka kvinnors deltagande , på ett sådant sätt att 40 procent av dem som får marie curie-stipendier , deltar i de rådgivande församlingarna och utvärderingspanelerna för hela det femte fou-ramprogrammet skall vara kvinnor .
för det ändamålet krävs en stimulans av debatten och erfarenhetsutbytet mellan medlemsstaterna , en samordningsstruktur för inrättandet av ett övervakningssystem inom det femte ramprogrammet , kallat &quot; kvinnor och vetenskap &quot; , vilket bl.a. skall sörja för insamling och spridning av statistik som samlats in under genomförandet av det femte ramprogrammet och som visar hur stor andel kvinnor som har deltagit i forskningsaktiviteterna .
i likhet med föredraganden anser jag att det fordras studier för att analysera orsakerna till skillnaden mellan det antal kvinnor som tar en naturvetenskaplig examen och det antal kvinnor som lyckas få en anställning på det området .
en bättre analys av de hinder som kvinnor stöter på gör att vi kan utveckla en strategi för att undanröja dessa hinder .
vi måste mobilisera de många nätverken med kvinnliga forskare och få deras hjälp för att formulera en gemensam forskningspolitik .
europaparlamentet kommer även i fortsättningen att uppmärksamt följa genomförandet av det femte ramprogrammet för fou , när det gäller främjandet av kvinnor , samt utformningen av idéer till riktlinjer för det femte ramprogrammet .
i fråga om vetenskap , forskning och europeiska unionens alla övriga politikområden , bör vi integrera genusdimensionen för att sätta stopp för den strukturella diskriminering som hindrar kvinnorna från att konkurrera med lika förutsättningar på arbetsmarknaden .
. ( fr ) i sitt meddelande om &quot; kvinnor och vetenskap &quot; framför europeiska kommissionen sina goda avsikter att berika den europeiska forskningen genom att mobilisera kvinnorna .
det är mycket bra och vi gläder oss åt det .
det finns faktiskt alltför få kvinnor som deltar i forskningsarbeten inom europeiska unionen .
vi vet att det enda vi kan göra för att förändra denna situation med underrepresentation av kvinnor inom det vetenskapliga området är att utveckla en utbildningspolitisk inriktning som systematiskt uppmuntrar en diversifiering av unga flickors yrkesval , och då de tagit sin examen vidta positiva åtgärder i arbetslivet .
men uppenbarligen har vissa kolleger tagit till brösttoner , med tanke på en punkt i betänkandet från utskottet för kvinnors rättigheter och jämställdhetsfrågor som bidrar till förvirring . en del tolkar den som en kvot , vilken skulle kräva 40 procent kvinnor inom den europeiska forskningen .
men så förhåller det sig givetvis inte , eftersom en sådan kvot skulle vara orealistisk .
i betänkandet nämns för övrigt inte när en sådan kvot är tänkt att uppnås .
för att skapa lugn och försäkra kollegerna har jag ingivit ett ändringsförslag till resolutionen , där vi helt enkelt noterar att kommissionen i sitt meddelande åtar sig att göra stora insatser för att öka kvinnors deltagande i gemenskapens forskningsprogram , vilket trots allt är hedervärt .
och varför inte notera att kommissionen skriftligen har meddelat att den anser 40 procent vara ett mycket viktigt mål för kvinnors deltagande på alla nivåer i genomförandet och förvaltningen av forskningsprogrammen .
detta är inte en kvot !
det är en mycket välgrundad avsiktsförklaring från kommissionens sida , i den mån det gäller dess egna och inte medlemsstaternas program .
staterna borde dock komma på den goda idén att för en gångs skull följa kommissionens goda exempel och sätta in lika stora insatser inom ramen för sina egna forskningsprogram .
men förutsättningen är givetvis att man inser det !
. ( fr ) det är lyckosamt att det fanns ett så stort samförstånd i debatten om mcnallys betänkande , som syftar till att utöka och underlätta kvinnors deltagande i yrken inom området för forskning och vetenskap .
i den här frågan vore det önskvärt att begreppet lika möjligheter får ett bättre genomslag i vardagen , och jag kan endast glädjas åt genomförandet av en politik som bidrar till att kvinnors legitima strävanden tillmötesgås : att få lika tillträde till vetenskapliga studier , att nå ansvarsposter som verkligen står i relation till deras resultat och förmåga , att se snabbt genomförda följdåtgärder som gör att de kan förena familje- och yrkeslivet .
detta är en nödvändig realistisk och pragmatisk politik , vars syfte är att avskaffa konkreta hinder som har konstaterats vara obestridliga orsaker till denna ojämlikhet . men enligt vår mening måste den absolut ta avstamp i begreppet komplementaritet , vilket är det enda som kan rättfärdiga en viljestark politik i frågan .
det är genom att respektera dessa värden , som verkligen innefattar en respekt för skillnader , och inte genom att luta sig mot ett påstående om en jämlikhet mellan könen - som i sig bär på motsägelser - som vårt reflektionsarbete och åtgärder måste koncentreras på i framtiden .
det finns i alla fall ingenting som motiverar att man gör det enkelt för sig och bedriver en kvantitativ politik , dvs. att införa kvoter . det skulle strida mot det medborgarskapsbegrepp som ledamöterna i uen-gruppen är särskilt måna om , och det skulle förmodligen få konsekvenser som står i motsats till dem som tycks eftersträvas i mcnallybetänkandet , nämligen att kvinnor skall delta i yrken på området för vetenskap och forskning i proportion till deras värde .
genom att kvinnorna får tillfälle att uppvisa sina verkliga förtjänster och så långt det är möjligt undanröja de hinder som är förknippade med deras särskilda villkor - dock inte inom ramen för en konflikt där de ger intryck av att angripa männens privilegier - kommer de att bevisa intresset av att underlätta utvecklingen av sina yrkeskarriärer , och därmed kommer de att uppnå en förändring av den balans som alltför ofta är till deras nackdel .
eftersom europaparlamentet har valt att rösta för en text som uttryckligen vädjar om en kvoteringspolitik , något som jag med stor beslutsamhet försökte kritisera i mitt yttrande , och trots att jag till stor del instämmer i de allmänna riktlinjerna , var jag tvungen att avstå från att rösta om betänkandet av mcnally .
andrabehandlingsrekommendation ( a5-0006 / 2000 ) av florenz
fru talman , ärade damer och herrar , kära kolleger ! vi har i dag i en andra behandling röstat om ändringsförslagen till direktivet om uttjänta fordon .
jag röstade emot hela direktivet , även på grund av att ändringsförslag 34 till artikel 12 och ändringsförslagen till artikel 5.4 inte fann tillräcklig majoritet här i kammaren .
jag kommer från ett land där 50 procent av eu : s bilpark tillverkas , och det är just det kostnadsfria återtagandet av det gamla bilbeståndet som är kostnadsintensivt och oacceptabelt .
här kommer enligt min åsikt även arbetsmarknaden att belastas väsentligt genom de kostnader som dessa företag kan vänta .
detta kan inte vara bra i en europeisk union där vi dagligen funderar kring sysselsättning .
jag anser att detta är en graverande brist som i princip inte heller passar vårt rättssystem .
ur denna synvinkel anser jag inte att detta direktiv är godtagbart .
fru talman ! jag skulle vilja yttra mig om florenz betänkande .
jag tycker att omröstningen har visat att rådets gemensamma ståndpunkt har försvagats men att de stora grupperna här - i synnerhet de tyska företrädarna för de stora grupperna - tack och lov inte lyckades förstöra själva kärnan i direktivet , nämligen producentansvaret .
tyvärr fick det passera att en effektiv ekologisk politik för avfallsströmmar nu försvagas , nämligen genom den obligatoriska riskbedömningen av ämnen vars hälsovådliga effekter egentligen har varit kända i flera år .
vi vet att bly , kvicksilver , kadmium och sexvärt krom gömmer stora toxiska faror och hälsorisker och att man genom talrika gemenskapsdirektiv har lyckats minska användningen av detta utan att det har förelegat någon riskanalys .
här har europaparlamentet tyvärr böjt sig för industrins intressen .
jag är likväl mycket glad över att man har inte har lyckats få majoritet för ändringsförslagen från florenz , lange och andra , vilka verkligen har försökt baxa ut producentansvaret och överlåta helt åt konsumenterna att stå för kostnaderna för en miljöanpassad hantering av uttjänta fordon .
jag tycker att det var ett försök som man verkligen borde skämmas över , och jag är glad att det inte lyckades , att man här inte lyckades samla majoritet för det som en stor regering och ledamöterna från en stor medlemsstat försökte sig på , nämligen att på grundval av deras nationella industris intressen dominera europaparlamentets hållning vid omröstningen .
fru talman ! trots att jag tillbringat större delen av mitt liv i snabba bilar håller jag med min kollega florenz om att man i direktivet om uttjänta fordon måste klargöra att direktivet inte omfattar veteranbilar .
dessa fina bilar är inte något avfall .
det var därför jag röstade för ändringsförslagen .
veteranbilarnas ålder skall inte heller fastställas eftersom det är stora skillnader mellan de nationella bestämmelserna .
på det här sättet kan man bevara historiskt värdefulla fordon för kommande generationer .
vi får inte heller glömma dem som har veteranbilar som hobby , deras antal överstiger 50 000 bara i finland .
i stillhet utför de ett mycket värdefullt kulturhistoriskt arbete .
. processen i parlamentet rörande denna fråga har varit minst sagt förvirrande .
inför omröstningen i plenum har nya ändringsförslag lagts fram , sådana som redan röstats ned i utskottet .
i den splittrade situation som nu uppstått anser vi därför att rådets skrivningar är de bästa .
vi behöver ett direktiv på detta område , och därför vill vi också undvika en komplicerad förlikningsprocess .
direktivet om uttjänta fordon kommer att statuera exempel för kommande lagstiftning .
det är därför viktigt att producentansvaret är tydligt ; det får inte på något sätt äventyras .
i dag granskar parlamentet för sista gången denna text om så kallade uttjänta fordon och deras öde , dvs. förstörelsen av dem , vilket är en lovvärd avsikt med respekt för vår miljö .
men det finns två aspekter som man absolut bör beakta i texten .
först och främst det finansiella ansvaret för denna förstörelse .
låt oss se till att det inte alltid blir densamme som betalar , dvs. fordonsägaren .
denne är redan tillräckligt beskattad för sitt fordon som i finansiellt hänseende inte är annat än en bottenlös källa .
helt nyligen har vi kunnat tala om principen att den som förorenar skall betala , låt oss då tillämpa den förnuftigt och med eftertänksamhet , utan ideologi och utan att ta miste på mål .
den andra grundläggande punkt som bör återfinnas i denna text , är en uttrycklig föreskrift om att samlarfordon inte skall omfattas av tillämpningsområdet .
på sina håll sägs det att man inte behöver skriva det , eftersom det är uppenbart , men jag är angelägen om att det görs , för vi har allt intresse av att anta tydliga texter .
låt oss därför rösta igenom dessa ändringsförslag för att bevara bilindustrins juveler .
dessa antika fordon bär vittne om en kultur och en passion som bör erkännas och respekteras av europa , i annat fall riskerar vår specifika karaktär att urvattnas .
det saknas inte exempel bland eu-texterna - i det fallet vet vi att luddighet eller oklarhet inte sällan leder till betydande tvister eller debatter .
jag skall bara nämna direktiven 79 / 409 och 92 / 43 .
tydliga texter är en garanti och en rättslig säkerhet för dem som dagligen kommer att tillämpa eller omfattas av dessa texter .
parlamentsledamöternas kallelse är inte att skapa tvister eller förse domare med rättegångsprocesser , vilka de än är , för då skulle vi inte uppfylla vårt uppdrag .
vi parlamentariker bör tvärtom anta kristallklara texter för att begränsa tvister .
( nl ) att florenzbetänkandet har gjort så mycket väsen av sig bevisades av den starka lobbymaskin som sattes in , såväl av industrin som av miljörörelsen .
jag beklagar att konstruktörerna bombarderade europaparlamentet och rådet med en hel rad argument som antingen inte höll eller som var falska .
jag vågar säga detta eftersom jag gjorde mig besväret att också ge mig ut på fältet och inhämta upplysningar hos bland annat skrotningsföretag som redan ägnar sig åt återvinning av bildelar med framgång .
de gjorde klart för mig att argumenten om till exempel säkerhetsrisker är struntprat .
billobbyn lyckades inte i dag , och det är jag glad för .
direktivet står fortfarande kvar .
jag räknar med att vi under förlikningen kommer att uppnå ett utmärkt resultat och att ansträngningarna för en bättre miljö vinner över orimliga industriella krav .
. ( en ) mitt parti har motsatt sig denna åtgärd och de föreslagna ändringsförslagen .
det finns få saker som är så säkra i livet som skatter , död och miljöförstörelse .
men det finns inte heller något som är så säkert som att eg : s miljödirektiv har lovvärda syften men i själva verket misslyckas med att uppnå fastställda mål .
när det gäller miljöförstöring liksom synd är vi alla emot den , men för den sakens skull får vi inte tro att varje åtgärd som föreslås mot detta onda med nödvändighet är god .
faktum är att detta direktiv , liksom så många andra som behandlar miljöfrågor , inte är bra .
som så ofta är fallet tillför det bara ännu en tung byråkratisk struktur för att kontrollera ett problem , vilket bara tjänar till att skapa flera arbetstillfällen för tjänstemän och kostar motorindustrin och konsumenterna en hel del pengar .
det enda det inte kommer att göra är att lösa problemet - det är att skjuta myggor med kanoner .
ingen , inte minst mitt parti , kan vara av någon annan åsikt än att återvinning skall främjas , men det bästa sättet att uppnå detta är att arbeta med marknaden , inte att skapa ett nytt byråkratiskt missfoster .
ett lämpligare sätt att gynna återvinning är sålunda att lägga skatt på producenter som inte ökar mängden återanvändningsbart material i sina fordon , detta för att med hjälp av skatteincitament och hjälp att rätta sig efter miljökrav uppmuntra privata återvinningsföretag samt skapa incitament för användning av återvunnet material .
självklart är detta områden där eu inte har någon jurisdiktion och inte heller skall ha någon sådan jurisdiktion .
i avsaknaden av sådan makt , borde man likväl inte försöka ersätta detta med en mindre effektiv åtgärd .
i stället borde man låta medlemsländerna utveckla sina egna system och undvika tendensen att ingripa där detta inte är önskvärt eller gör någon nytta .
betänkande ( a5-0007 / 2000 ) av berger
med detta förslag till direktiv vill man fastställa villkoren för utstationering av arbetstagare från tredje land i samband med tillhandahållande av tjänster över gränserna .
nationaliteter från tredje land med legalt uppehållstillstånd i en medlemsstat åtnjuter inte rätten till fri rörlighet i europeiska unionen .
hittills har det varit stränga restriktioner i den fria rörligheten för arbetstagare från länder utanför unionen .
det är alltså positivt att man underlättar rörligheten för arbetstagarna i europeiska unionen , även för arbetstagare från tredje land .
emellertid syftar bara diektivförslaget till att tillåta deras förflyttning till en annan medlemsstat när det är i arbetsgivarens regi , en arbetsgivare som är etablerad i ett land där han också har sin hemvist , men möjligheteten till rörlighet är begränsad till tiden för utstationering , och bara till den medlemsstat där arbetstagaren har blivit utstationerad .
detta innebär att det främsta syftet med detta förslag inte är att lösa problemet med dessa arbetstagares rörlighet , utan bara att skapa bättre villkor för företagen som tillhandahåller tjänster .
å andra sidan för att underlätta förfarandena tas det i bergerbetänkandet upp ändringsförslag som är djupt diskutabla , vilket skapandet av ett gemensamt informationssystem om tillgång till kort eg-kort utgivna av en myndighet i någon av medlemsstaterna är ett exempel på .
betänkande ( a5-0007 / 2000 ) och ( a5-0012 / 2000 ) av berger
. ( fr ) det är med största tillfredsställelse som jag välkomnar de två förslag till direktiv som syftar till att underlätta den fria rörligheten för arbetstagare från tredje land och samtidigt det fria tillhandahållandet av tjänster .
dessa förslag går i huvudsak ut på att införa ett eg-kort för tillhandahållande av tjänster , som i framtiden kommer att ge nära 5 miljoner medborgare från tredje land som vistas legalt i en av europeiska unionens medlemsstater möjlighet att tillhandahålla tjänster i andra medlemsstater , något som i dag hindras av problem med att få visum och arbetstillstånd .
det första förslaget i direktivet skall tillåta de företag som är etablerade i en medlemsstat och som har arbetstagare från tredje land att tillfälligt utstationera dessa arbetstagare i en annan medlemsstat för att tillhandahålla tjänster där .
i enlighet med de föreskrivna bestämmelserna skall arbetsgivaren bara behöva göra en förfrågan om ett kort för tillhandahållande av tjänster för varje berörd arbetstagare .
för att kunna få ett sådant kort bör arbetstagaren logiskt sett vistas legalt i en medlemsstat och omfattas av ett socialförsäkringssystem .
det andra förslaget ger samma rättigheter åt egna företagare från tredje land .
innehållsmässigt ansluter jag mig till europeiska kommissionens förslag .
vissa bestämmelser kan dock skapa förvirring , och därför röstar jag för de ändringsförslag som har ingivits av föredraganden .
de kan bidra till att bestämmelserna tydliggörs och således till att man förekommer alla former av missbruk !
andra ändringsförslag syftar till att förenkla de administrativa förfarandena , till exempel genom att låta medlemsstaterna utse en myndighet som skall ha ansvaret att utfärda korten .
en sådan ändring verkar nödvändig för att undvika det byråkratiska krångel som alltför ofta bromsar en bra tillämpning av nya bestämmelser .
därför kan jag bara glädja mig åt att dessa ändrade direktiv har antagits , eftersom vi inte mycket längre kan acceptera att personer som under lång tid har vistats legalt inom europeiska unionen skall stöta på så många svårigheter .
det går stick i stäv med den grundläggande princip om icke-diskriminering som är inskriven i unionens grundfördrag .
betänkande ( a5-0003 / 2000 ) av marinho
. den stundande regeringskonferensens viktigaste uppgift är att reformera eu inför mottagandet av de nya medlemsländerna .
vi stöder därför givetvis att europaparlamentet nu ger sitt formella klartecken till att regeringskonferensen startar .
vi anser dock att regeringskonferensen skall begränsas till frågor som är nödvändiga för att utvidgningen skall kunna göras .
detta hävdade vi också i november 1999 , och vi vill därför hänvisa till vår röstförklaring av den 18 november 1999 .
( fr ) i den ståndpunkt som europaparlamentet just har antagit om inledningen av nästa regeringskonferens , vädjar parlamentet om att man bör &quot; inleda en konstitutionell process &quot; .
denna vilja att kontrollera nationerna med en juridiskt sett högre stående text kommer också till uttryck på de första sammanträdena i den församling som har i uppdrag att utarbeta en så kallad stadga om de grundläggande rättigheterna , men i realiteten en maskerad konstitution .
den viljan uttrycks också i det osannolika steg som i dag tas i europaparlamentet : önskan att radera resultatet av de fria valen i österrike genom att rösta igenom en resolution .
samma vilja att göra nationerna till vilka underordnade administrativa regioner som helst , framgår också av alla sidorna i kommissionens yttrande inför regeringskonferensen .
den centrala idén består i att generalisera omröstningarna med kvalificerad majoritet och samtidigt förändra innebörden av denna kvalificerade majoritet , genom att omvandla den till en dubbel enkelmajoritet - staterna och befolkningarna - med syftet att öka kommissionens handlingsutrymme och minska densamma för de stater som är i minoritet .
fransmännen kommer utan tvekan att vara intresserade av att - så här i förbigående - få veta att kommissionen begär en ändring av artikel 67 i amsterdamfördraget för att där införa majoritetsomröstningar , samt ett medbeslutande med europaparlamentet .
man bör minnas att denna artikel , som handlar om invandringspolitikens överföring till gemenskapspelaren , föreskriver att besluten skall fattas enhälligt i rådet under fem års tid , och att rådet sedan skall bedöma om det eventuellt är lämpligt att ändra på systemet .
i frankrike , både i nationalförsamlingen och i senaten , kände sig många parlamentsledamöter lugnade när fördraget ratificerades , eftersom man sade att rådet under alla omständigheter kommer att ha frihet att välja och att det därmed skulle kunna bevara enhälligheten .
men i dag föreslår barnier - den europaminister som förberedde amsterdamfördraget och som under tiden har blivit ledamot av europeiska kommissionen - att man vid nästa regeringskonferens skall besluta att rådet skall arbeta på de här frågorna med majoritetsbeslut .
detta är ett exempel på att vi ständigt hamnar i en ond cirkel när vi spelar spelet om den europeiska integration med institutionerna i bryssel .
fransmännen måste inse att alla dessa åtgärder inte endast syftar till att deras land skall försvinna såsom ansvarigt beslutscentrum , utan att man också kommer att utnyttja alla medel för att avtvinga dem deras samtycke till detta .
ger de efter är de förlorade .
för det man håller på att ta bort , det är deras försvarsmedel , ett efter ett .
( da ) de danska socialdemokraterna har i dag röstat emot betänkandet om sammankallande av regeringskonferensen .
det är avgörande för oss att denna regeringskonferens kan avslutas före utgången av år 2000 , så att det inte blir formella förhållanden som röstviktning i ministerrådet och sammansättningen av kommissionen och europaparlamentet som lägger hinder i vägen för utvidgningen av eu .
vi var därför också mycket nöjda med de beslut som fattades om detta på toppmötet i helsingfors i december .
en alltför ambitiös utvidgning av dagordningen vid nuvarande tidpunkt riskerar att försena utvidgningsprocessen .
detta vill vi inte skall ske - vi har därför röstat emot .
vi håller emellertid helt med våra kolleger om att det finns behov av öppenhet i samband med regeringskonferensen , så att medborgarna får klart för sig hur arbetet fortskrider .
vi är nöjda med att det sattes upp en begränsad dagordning för regeringskonferensen vid mötet i helsingfors .
utformningen av det framtida eu bör även eventuella blivande medlemsstater vara med och ha ett inflytande över .
valet till europaparlamentet 1999 visade med all tydlighet att medborgarna inte följer med i tankegångarna om ett allt mer brysselfederalistiskt eu .
. ( fr ) när nästa regeringskonferens inleds blir europeiska unionens metod åter aktuell .
än en gång kommer stats- och regeringscheferna att skaffa sig ensamrätt till debatten .
det betyder att femton personer kommer att diskutera och fatta beslut inom lykta dörrar om 350 miljoner människors framtid .
man kan därför förstå folkens ointresse för ett europeiskt bygge som uppförs bakom ryggen på dem och långt ifrån deras angelägenheter .
det räcker faktiskt med att titta på regeringskonferensens dagordning : institutionerna , utvidgningen och ett självständigt försvar .
i realiteten handlar det om att förstärka den verkställande makten , att utveckla östländernas införlivande av liberalismen och att driva på en militarisering av europa , bl.a. genom att utöka försvarsbudgetarna .
det sociala europa , något som eu framhåller , har helt enkelt försvunnit från dagordningen .
allt detta legitimerar bara utvecklingen av motståndsrörelser på europanivå , rörelser som vill införa en social stadga för att arbetstagarnas viktigaste krav skall harmoniseras ovanifrån .
jag röstade för resolutionen som är positivt till sammankallandet av en regeringskonferens eftersom det befäster det portugisiska ordförandeskapets filosofi , med stöd från en stor majoritet i parlamentet , om att öppna regeringskonferensens dagordning för andra frågor än de som är strikt relaterade till maktbalansen mellan medlemsstaterna , stora och små , så som ursprungligen fastställdes i kallelsen till rådet i helsingfors .
tyvärr är de ämnen som tas upp i resolutionerna om de framtida frågorna för en revidering av fördraget om behovet att se över artikel 7 , som handlar om avstängning av en medlemsstat om den på ett allvarligt och återkommande sätt kränker unionens ursprungliga principer i artikel 6 .
så som visas i den nuvarande krisen med österrike , har unionen rätt att försvara sig .
emellertid är de rättsliga mekanismerna som finns i fördraget svaga , och svåra att tillämpa politiskt och rättsligt , de klassificerar inte institutionernas makt och garanterar inte en rättslig behandling av en process av större betydelse vilket just ett fördömande och avstängning av en medlemsstat innebär .
därför anser jag att denna fråga genast måste föras upp på regeringskonferensens dagordning , och detta motiverar i sig en långtgående revidering .
de frågor , som vi för närvarande anser vara centrala , när det gäller sammankallande av en regeringskonferens för att revidera fördragen är långt viktigare än kontroversen här angående varje dagordnings dimension , när det gäller möjligheten att formulera förslag till nya frågor att ta upp och europaparlamentets deltagande i den .
de relevanta frågorna , enligt vår mening , handlar om regeringskonferensens möjligheter och syften och de frågor som kommer att debatteras .
vi tvivlar på möjligheterna eftersom vi har de verkliga målen i sikte , kanske långt ifrån det alltid nämnda anpassningen till den planerade utvidgningen .
detta syns särskilt i det innehåll som eftersträvas , speciellt inom de områden som ej löstes i amsterdam - och detta tyder på ett framtida skapande av oacceptabla direktorat - , men också för det som handlar om andra och tredje pelaren , vilka tenderar i en riktning mot en oönskad militarisering av europeiska unionen .
det här är några av de främsta skälen till att vi inte stöder inriktningen av detta resolutionsförslag .
. för att kunna påverka utvecklingen måste europaparlamentet inta en mer konstruktiv attityd till regeringskonferensens dagordning än som framkommer i denna resolution , vilken i alltför stor utsträckning ägnar sig åt besvikelse och negativism över det beslut som europeiska rådet fattade i helsingfors i december 1999 .
europaparlamentet och dess konstitutionella utskott borde i stället ha preciserat sig och koncentrerat sig på några få punkter utöver rådsbeslutet i helsingfors och därmed ange vad man anser vara mest angeläget att ta upp till behandling , bland annat frågan om inrättande av en åklagare för brottslighet riktad mot europeiska unionens institutioner och deras ekonomiska intressen .
vi svenska kristdemokrater motsätter oss också hot om att försena östutvidgningen av eu som framförts om inte regeringskonferensen utvidgas mycket omfattande utöver vad som blev kvar från förra regeringskonferensen i amsterdam 1997 .
- den stundande regeringskonferensens viktigaste uppgift är att reformera eu inför mottagandet av de nya medlemsländerna .
jag stöder därför givetvis att europaparlamentet nu ger sitt formella klartecken till att regeringskonferensen startar .
jag anser dock att regeringskonferensen skall begränsas till frågor som är nödvändiga för att utvidgningen skall kunna genomföras .
i övrigt hänvisar jag till min röstförklaring av den 18 november 1999 där jag klargör min inställning gentemot överstatlighet och ett gemensamt försvar .
gemensam resolution om österrike
fru talman ! gruppen nationernas europa har inte anslutit sig till ppe-de- och pse-gruppens gemensamma resolution om den politiska situationen i österrike , vilken uppstått till följd av att de konservativa och jörg haiders nationalliberaler bildat koalitionsregering .
ppe-de- och pse-gruppens resolution applåderar det initiativ som togs av fjorton medlemsstater för att sätta press på österrike , genom att organisera en sorts diplomatisk bojkott .
det som chockerar oss mest är att denna gemensamma intervention viftar med fördragets principer som om det någonstans stod skrivet att ett folks fria och demokratiska uttryck kan upphävas av grannländernas stats- och regeringschefer , som för övrigt har aktat sig noga för att samråda med sina respektive folk .
vilka verbala övertramp jörg haider än har gjort , och vi beklagar faktiskt dem , har österrikarna gjort ett demokratiskt val , och det måste vi respektera .
i våra ögon är det uppenbart att vänstern i europaparlamentet - i samförstånd med den österrikiska vänster som besegrades i striden om väljarna - har iscensatt en ren och skär politisk operation som för tankarna till en olycksbådande epok , men som vi lyckligtvis har lämnat bekom oss .
även om jämförelsen mellan haider och hitler saknar all trovärdighet , har den delvis fyllt sin funktion genom att få vissa ppe-de-ledamöter att vackla .
men bortsett från denna politiskt förslagna operation , finns det en sak som majoriteten i europaparlamentet särskilt fruktar , och det är att ifrågasättandet av vänsterns och högerns sammanboende i österrike - något som har fördärvat det politiska livet - snart sprider sig till det europeiska systemet med gemensamt styre , ett styre som ger upphov till lika beklagansvärda effekter .
för att undvika ett sådant ifrågasättande är denna majoritet beredd till allt : att sudda ut resultaten av fria val ; att inrätta en tankepolis ; att införa en ny form av totalitarism .
fru talman ! för ledamöterna från nationella fronten , vlaams blok och den italienska sociala rörelsen vill jag ställa följande fråga : vem är det som drar i trådarna i den förskräckande inblandning i österrikes inre angelägenheter som europeiska unionen har hängett sig åt i strid med den allmänna internationella rätten , i strid med fördragen , i strid med moralen ?
är hysterin spontan ?
är den en frukt av ren dumhet eller - mera troligt - av en avsiktlig strategi , densamma som brukas överallt annars i världen ?
vem dikterar sin vilja för de europeiska nationerna och gör anspråk på att förbjuda dem att välja ett eget öde ?
hemliga nätverk ?
regeringen i washington ? den i israel ?
eller deras socialistiska reservtrupper , som i denna församling har fräckheten att sprida sina värderingar bland oss ?
vilka är då socialisternas värderingar , de socialister som har nått stora valframgångar under det senaste seklet genom att förespegla de sämst lottade en större social rättvisa , men som i dag inte är mer än ett parti för skyddade tjänstemän , etablerade fackföreningar och statskapitalism ?
vilka är det belgiska socialistpartiets värderingar , ett parti som går från pedofilskandaler till korruptionsaffärer , till att börja med vandamaffärerna , såsom agustaaffären ?
vilka är värderingarna inom det franska socialistpartiet , som i urba- , sages- och graco-affärerna har övat utpressning mot alla de kommuner som är beroende av socialisterna ?
i françois mitterrands parti , mitterrand som tilldelades vichyregimens emblem av pétain , har de högsta ämbetsmännen just blivit tagna på bar gärning , när de levde gott på att förskingra offentliga medel avsedda till en sjukförsäkring för studenter .
jag skall inte ta upp det italienska socialistpartiets korruptionsaffärer , för man slår inte på den som redan ligger , och än mindre på den som redan är död .
jag skall däremot tala om det spanska socialistpartiet , som just har ingått en allians med slaktarna från albacète som gjorde upp med de baskiska nationalisterna med hjälp av lejda mördare .
jag kommer att tala om det tyska socialistpartiet , som har för avsikt att undervisa oss om andra världskriget - ett international-socialistiskt parti , precis som dess likar var national-socialistiska , som fortfarande marscherar , waffen-ss : s parti ...
fru talman ! jag har haft stora svårigheter med denna resolution .
till slut lade jag av flera orsaker ned min röst .
jag sympatiserade med edd-gruppens ändringsförslag , som behandlar förkastandet att eu : s ingriper i bildandet av regeringar i medlemsstaterna , men jag var tvungen att lägga ned min röst , eftersom förslaget precis följde på fördömandet av främlingsfientlighet , rasism etc. och jag tyckte att det kunde misstolkas .
men jag funderar över hur klokt detta är .
för det första uppstår frågan om bekämpning av intolerans med intolerans och de långsiktiga följderna av detta .
jag undrar också hur klokt det är av eu att reagera på regeringsbildningen i österrike och hur detta kommer att påverka den allmänna opinionen där .
för tillfället verkar det som om haiders parti snarare får mera stöd än mindre från oppositionen i utomstående regeringar .
till och med usa har nu meddelat att man överväger att bryta de diplomatiska förbindelserna .
vi undrar om detta inte i själva verket underblåser främlingsfientligheten och gagnar de partier och människor som understöder detta .
jag tycker verkligen att folk borde vara väldigt försiktiga .
om man vill bekämpa främlingsfientlighet och rasism , och jag tror att vi måste det , måste vi fokusera på grundorsakerna .
vi måste iaktta de människor som röstar på dessa partier och förstå varför denna situation uppstår .
det är ingen situation som de flesta i detta parlament önskar , men vi måste vara försiktiga i vårt val av synsätt , så att vi inte till slut åstadkommer raka motsatsen till det vi försöker uppnå .
fru talman , kära kolleger ! jag avvisar varje sorts främlingsfientliga och rasistiska uttalanden , manifestationer eller känslor .
jag försvarar intensivt de mänskliga rättigheterna och rättsstaten , vilket europa består av .
men jag är ändå oense med det befängda agerandet som ordförandeskapet ( tyvärr det portugisiska ordförandeskapet ) har initierat i en verkligt institutionell dumhet för fjorton andra medlemsstaters räkning .
detta är inte ett sätt att bekämpa extremism på .
det kan till och med vara ett sätt att spela dem i händerna på ett oöverskådligt sätt .
den kaskad av förvirrade och förhastade åtgärder som vräkts över österrike blandar ihop allt på ett oproportionerligt sätt , och det stör många medborgare med god vilja och utgör risker som inte har beaktats .
det finns en oförenlig motsättning mellan ståndpunkter som tas i de mänskliga rättigheternas och rättsstatens namn , men som , samtidigt förolämpar österrikarna i grundläggande rättigheter och kör över de grundläggande rättigheterna i en rättsstat , i detta fall fördragets bestämmelser .
vad vill vi när vi inleder en regeringskonferens ?
ett europa med 27 länder eller ett europa med 14 , eller ännu mindre ?
vi är för europa , ett europa som hedrar alla de steg vi har tagit för att komma hit , ett europa som respekterar fördragen och lagen , ett europa där österrike behövs .
det är viktigt att säga detta !
fru talman ! jag är glad och stolt över att detta parlament , med övervägande majoritet , har fördömt bildandet av koalitionen i österrike med haiders liberala parti .
haider har under de senaste åren såväl i ord som handling visat att han förtjänar att utestängas från en vanlig demokratisk dialog .
han har inte bara beundrat adolf hitler , berömt waffen ss och vägrat fördöma en terroristattack som dödade fyra romer , han har också varit ledamot i det regionala styret i kärnten .
han har lett satsningar för att dra in bidrag åt österrikes slovenska minoritet och stöd åt immigranter .
en del har hävdat att vi inte har rätt att ingripa i österrikisk politik .
de har fel .
genom europeiska unionens fördrag är vi förpliktade att skydda grundläggande rättigheter .
en del har hävdat att vi måste acceptera resultaten av demokratiska val .
men demokratiska val gör inte demokrater av dem som har hotat demokratin .
för dem som hävdade samma sak med avseende på tyskland under 1930-talet , finns det ett tragiskt minnesmärke i form av förintelsen - 6 miljoner judars död .
men vi skall inte döma haider för hans ambition .
somliga människor ändrar aldrig åsikt .
de skyldiga är egentligen kristdemokraterna i österrike som beter sig som syndabockar för att återuppliva det hot mot europa som vi trodde dog i berlin 1945 .
vi har nyligen antagit en resolution som fördömer jörg haiders liberala partis rasistiska och främlingsfientliga förflutna i österrike . detta har gjort det möjligt för våra regeringar att handla genom att bryta de politiska förbindelserna med varje regering som han är medlem i och visar också vårt stöd för anti-rasistiska grupper inom den demokratiska majoriteten av österrikes folk .
vi varnar för att den här koalitionen , om den bildas i dag , på ett oacceptabelt sätt legitimerar extremhögern , i direkt motsats till de principer om fred och försoning som för oss samman i denna europeiska union .
detta är de värderingar vi önskar se hos dem som vill gå samman med oss .
europaparlamentet kräver att europeiska kommissionen är vaksam när det gäller rasistiska aktioner i österrike och hotar med att utesluta österrike som medlem ur europeiska unionen om sådana förekommer .
jag är stolt över att understödja en sådan resolution .
trots att vårt förslag om att dra tillbaka alla politiska inbjudningar till österrikiska regeringsföreträdare till europaparlamentet inte antagits i dag , vill jag meddela att vi kommer att fortsätta med att driva detta förslag för att säkerställa att europaparlamentet gör allt som står i dess makt för att bekämpa återkomsten av nynazister till regeringar i europa .
jag respekterar parlamentets önskan som den har framkommit , men jag måste också säga att folkens rätt till självbestämmande inte kan ifrågasättas ens av europaparlamentet .
handlingen är orättvis gentemot våra österrikiska kolleger , både nationella och europeiska parlamentsledamöter , och luktar misstänksamhet och politiska , men också kommersiella , intressen lång väg .
jag tycker inte att man botar medborgarnas ointresse för europa med dessa signaler .
den österrikiska extremhögern har fått en oförtjänt present .
jag uppskattade de italienska radikalernas ståndpunkt mycket , och det säger jag utan att förglömma de historiska och faktiska skillnaderna mellan italienska och österrikiska liberaler .
jag har under många år i ord och handling varit engagerad i den antifascistiska kampen , kampen för jämställdhet och kampen mot främlingsfientlighet .
men det som skett under den senaste tiden , först i samband med det som i verkligheten var problem inom ministerrådet , sedan med ordförande prodis problem med den österrikiske kommissionären och senast i och med denna resolution , är inte något jag kan ställa upp på .
jag har inte kunnat rösta för denna resolution , även om jag stöder vissa slutsatser .
det handlar först och främst om en illavarslande blandning av makt , arrogans och svaghet från den europeiska unionens sida .
dessa åtgärder strider inte bara mot fördragen och ger unionens organ mer maktbefogenheter än vad som tillkommer dessa , utan det värsta är att de kommer att motverka sitt eget syfte .
det kommer inte att försvaga haider och fpö ( österrikiska liberala partiet ) , det kommer tvärtom att stärka dem .
vi uppnår det rakt motsatta .
på detta sätt bekämpar man inte rasism och högervridning .
( da ) venstres ledamöter vid europaparlamentet lägger vikt vid att parlamentet vid antagandet i dag inte har stött de fjorton statsministrarnas diplomatiska sanktioner mot österrike .
därför stödde venstres ledamöter vid parlamentet det liberala beslutets kraftfulla avståndstagande från varje form av främlingsfientlighet i österrike och på andra ställen .
vi fäster avgörande vikt vid att amsterdamfördragets nya bestämmelser används om detta är nödvändigt , så att ett land som i handling kränker grundläggande medborgerliga rättigheter genom diskriminering e.d. , fråntas rösträtten i eu : s ministerråd ( art . 7 ) .
. ( el ) fpö : s deltagande i österrikes regering innebär en mycket stor fara för europeiska unionens fortsatta politiska utveckling .
det rör sig om &quot; ormens ägg &quot; som nu tyvärr åter dyker upp i europa , starkare än någonsin sedan andra världskriget .
europaparlamentet och unionens regeringar är skyldiga att politiskt isolera en regering som innehåller anhängare av nazism och främlingsfientlighet .
europeiska unionen - och samtidigt de båda dominerande politiska riktningarna , socialdemokrater och kristdemokrater - har ett stort ansvar , för det är genom emu : s dogmatiska och stränga budgetpolitik , nedrustningen av välfärdsstaten och hyllandet av den tygellösa konkurrensen som stora befolkningsgrupper har marginaliserats , och därigenom har högerextremistiska demagoger av haiders typ fått möjlighet att mobilisera anhängare till sin nynazistiska politik .
( fr ) eftersom europaparlamentets bestämmelser inte tillåter oss att lägga fram en egen resolution för att fördöma haiders parti , liksom alla partier från vilket europeiskt land som helst som sprider rasistiska , främlingsfientliga och illvilliga tarvligheter mot invandrade arbetstagare , har vi röstat för kompromissresolutionen utan att stämma in i flera bedömningar och ordalag , för att visa vår solidaritet med dem i österrike som motsätter sig den österrikiska extremhögern och dess demagogi .
vår röst innebär på intet sätt en garant för de partier som undertecknat kompromissresolutionen , varken för deras nuvarande politik eller deras framtida attityd i händelse av ett ökat hot från extremhögern .
vissa av dessa partier , som ger sig ut för att vara republikanska och demokratiska , har anammat extremhögerns demagogi - av medbrottslighet eller valtaktiska skäl - om så bara för att - öppet eller på ett hycklande sätt - göra de invandrade arbetstagarna ansvariga för arbetslösheten och försvåra deras liv .
de personer från de undertecknande partierna som leder eller har lett en regering i europeiska unionens olika länder , har på ett mera allmänt plan en del av ansvaret för extremhögerns nyförvärvade inflytande , eftersom de bedriver en politik som av lojalitet med de stora arbetsgivarnas intressen saknar åtgärder för att bekämpa arbetslösheten och den misär som följer i dess fotspår , och därigenom underblåser extremhögerns främlingsfientliga demagogi .
. ( fr ) den här veckan har europa utan tvivel gett till sitt första politiska skrik .
genom att kraftfullt och snabbt fördöma det faktum att jörg haiders främlingsfientliga och antieuropeiska parti deltar i den österrikiska regeringen , vilket saknar motstycke sedan andra världskrigets slut , har europeiska unionen signerat sin politiska födelseakt och bekräftat att den inte endast är en ekonomisk och finansiell gemenskap , en stor marknad , &quot; affärsmännens europa &quot; .
just nu blottas en del av dess framtid , dess innersta väsen , dess själ .
för första gången har europaparlamentet kunnat göra sin röst hörd .
de europeiska socialdemokraternas upprop , på olivier duhamels initiativ , har väckt sinnena och möjliggjort ett beslutsamt och direkt politiskt gensvar på denna helt nya och oacceptabla situation .
14 europeiska stater har gett prov på denna beslutsamhet genom att enhälligt och omedelbart - med a. guterres röst - fördöma risken för en österrikisk politisk urspårning .
detta modiga ställningstagande inleder ett nytt kapitel i det europeiska byggets historia .
äntligen går vi tillbaka till ursprunget , en gemenskap uppbyggd på viljan att vända ryggen åt ett förflutet märkt av hat och utestängning och i stället ansluta oss till humanistiska värden som öppenhet och tolerans .
europa hade förmågan att resa på sig och fördöma det oacceptabla .
men med tanke på att det saknas juridiska instrument för denna politiska vilja - de sanktioner som föreskrivs i artikel 7 i fördraget är nästan omöjliga att tillämpa - kommer då europa att kunna hålla huvudet högt inför hotet om en systematisk blockering av hela den institutionella strukturen ?
i dag gäller det europas trovärdighet , innan vi i morgon kan ta emot de ännu sköra demokratierna i det f.d. östblocket .
europa måste nu omsätta sina ord i handling för att i allas ögon bekräfta hur stora våra återfunna ambitioner faktiskt är .
. ( fr ) när vi nu röstar om en gemensam resolution mot att nynazister skall ingå i en regering i europeiska unionen , måste jag beklaga att kompromisstexten framför allt saknar bestämdhet .
jag röstar för den , för det vore omöjligt att europaparlamentet inte skulle ta ställning efter gårdagens mycket utmärkta politiska debatt .
men personligen fortsätter jag att bekämpa extremhögern , jag fortsätter att samla in underskrifter till en petition för att kräva åtgärder som kan gå så långt som till att utesluta österrike och jag fortsätter genom att organisera en stor medborgardemonstration i lille på lördag kl. 15.00 .
fascismen och nynazismen är som cancer !
det djävulska djuret har väckts !
för mig är det inte tal om att låta dem utvecklas och frodas utan att slåss med stor energi .
europa föddes ur en vilja till fred , frihet och tolerans .
det kommer inte på fråga att europa skall acceptera att hysa främlingsfientliga , rasistiska och antisemitiska ministrar .
räkna inte med att jag förblir stum och passiv .
. ( en ) i gårdagens debatt i europaparlamentet uttryckte en del parlamentsledamöter oro över att vi lägger oss i ett medlemslands interna angelägenheter .
en sådan oro är onödig .
europaparlamentet har aldrig tvekat att kommentera en utveckling man inte samtycker till i medlemsstaterna .
vi har fördömt baskisk och irländsk terrorism .
vi har motsatt oss rasism och kränkningar av minoriteters rättigheter .
det är vårt ansvar som parlament , särskilt som europeiska unionens demokratiskt valda röst , att kritiskt kommentera den nuvarande politiska utvecklingen i österrike , vilken står i konflikt med parlamentets linje .
genom att kommentera och klargöra vår ståndpunkt hindrar vi inte något parti i österrike att bilda en koalitionsregering .
vi förklarar ändå för dem , vilket det är vår rättighet och plikt att göra , att ett sådant beslut , om de fortsätter på det sättet , kan leda till vissa konsekvenser och att vi i själva verket varnar dem på förhand .
andra påstår att vi borde skjuta upp domen tills vi ser detaljerna av en sådan överenskommelse .
ett sådant synsätt är inte bara en politisk smitning , det är uttryckligen farligt .
genom att nå en överenskommelse med jörg haider och hans parti , skulle de österrikiska kristdemokraterna i ett slag ge högerextremismen politisk legitimitet och dessutom ge dem tillgång till makt - vilket de kommer att använda som startplatta för ännu större valframgångar .
därför måste europeiska unionen klargöra sin ståndpunkt beträffande den nuvarande situationen i österrike .
. vi har röstat för den gemensamma resolutionen för att uttrycka vår solidaritet med alla dem som utsätts för främlingsfientlighet och rasism .
vi har också röstat för resolutionen i protest mot den avskyvärda politik jörg haider står för .
vi är dock mycket kritiska till de metoder de 14 medlemsländerna använt sig av i denna fråga .
i resolutionen saknas en tydlig hänvisning till respekten för medlemsländernas nationella identitet och konstitutionella traditioner i enlighet med artikel 6 i fördraget .
det saknas också en punkt om eu : s medansvar för den sociala och politiska utveckling i europa och österrike som varit en av förutsättningarna för haiders valframgång .
högerextremism är - idag , som tidigare i europas historia - resultatet av otrygga sociala och ekonomiska livsvillkor .
den nedskärningspolitik som följt i emu-anpassningens spår har befrämjat högerextremismens framgångar .
en radikal politik för trygghet och rättvisa i varje land är den bästa garantin för en demokratisk utveckling i europa .
denna förklaring avger jag på csu-gruppens vägnar .
det är outhärdligt att eu blandar sig i regeringsbildningen i en medlemsstat .
det tillkommer inte eu att göra så .
i stället för ett förhastat fördömande av fpö och den österrikiska regering som är under bildande fordras först och främst en kritisk undersökning och värdering av regeringsförklaringen och partiprogrammet samt koalitionens politik .
först efter att med kritiska ögon ha satt sig in i den kommande politik som de i koalitionssamtal inbegripna partierna ämnar driva har man möjlighet att avgöra huruvida denna regering strider mot europas demokratiska anda .
detta betyder inte att vi sympatiserar med haider .
csu : s europeiska parlamentsledamöter hyser inga som helst sympatier för fpö-ledaren haider .
som politiker måste vi tvärtom ställa oss frågan varför 27 procent av den österrikiska befolkningen valde ett parti som fpö vid valen i oktober 1999 .
vi måste analysera orsakerna till detta och försöka undanröja de orsaker som leder fram till sådana resultat .
endast en analys av fpö : s argument och politiska innehåll kan förhindra en radikalisering av politiken i österrike .
i europaparlamentets resolution frågar man däremot inte efter orsakerna till det österrikiska valresultatet och pekar heller inte på några möjliga lösningar .
detta är grunden till varför csu : s europagrupp uttalar sig mot resolutionen .
. ( fr ) &quot; ty han visste det som den jublande skaran var okunnig om och som man kan läsa om i böcker , nämligen att pestens bacill aldrig vare sig dör eller försvinner , att den under decennier kan slumra i möbler och källare , koffertar , näsdukar och pappersluntor och att den dag måhända skulle komma , då pesten , människorna till olycka och varnagel , ånyo skulle väcka sina råttor och sända dem ut att dö i en lycklig stad . &quot;
med dessa ord avslutar albert camus en lång allegorisk berättelse som beskriver oraninvånarnas svåra kamp mot pesten , för att efter andra världskrigets slut påminna oss om att kampen mot nazismen - &quot; den bruna pesten &quot; som den då kallades - inte kan krönas med en definitiv seger .
att rashatet , det främlingsfientliga våldet , rädslan och avvisandet av det annorlunda alltid kan återuppstå och komma att dominera vilken grupp av människor som helst , eftersom det är något som bottnar i människans lägsta sidor .
det är i denna bemärkelse de aktuella händelserna i österrike måste betraktas som tragiska .
för första gången sedan andra världskriget står ett öppet pronazistiskt , rasistiskt och främlingsfientligt parti på tröskeln till makten i ett europeiskt land .
inför detta hot - som i sig bär på ett förnekande av det europeiska byggets centrala idé - får ingenting stå i vägen : varken juridiska hårklyverier om vad fördraget tillåter och inte tillåter eller legitima frågetecken kring rätten till inblandning , eller en löjeväckande respekt för en formell demokrati , och framför allt inte den känsla av maktlöshet som griper oss inför en händelse som vi med våra övertygelsers fulla kraft vägrar att acceptera , men som vi inte har någon kontroll över .
som förtroendevald från ett franskt utomeuropeiskt departement , la réunion , en sammansmältningens och blandningens jordmån där befolkningen under de tre senaste seklerna har formats av successiva tillskott av européer , svarta från afrika och madagaskar , soldater från indien och pakistan och till och med kineser , upplever jag varje dag den djupaste sanningen i saint-exupérys ord : &quot; om du är olik mig , min bror , gör du mig inte illa , nej långt därifrån , du berikar mig ! &quot; .
det är den mänskliga mångfalden som har skapar vår främsta rikedom , och därför är det min plikt att förfölja och fördöma allt som kan kränka den - var den än visar sig .
av alla dessa skäl har jag med stor beslutsamhet röstat för den resolution om den österrikiska regeringsbildningen som lagts fram i kammaren .
. ( fr ) jörg haiders befordran , till följd av att fpö och den konservativa högern bildar regering , markerar en förfärande återuppståndelse av det monster som liberalismen skapat .
fpö : s framgångar har lika mycket att göra med de intyg om respektabilitet som tilldelats av den österrikiska högern och socialdemokratin som med de sistnämndas politik , vars sociala misslyckande har banat vägen för extremhögerns populism .
i resolutionen aviseras eventuella diplomatiska åtgärder för att politiskt isolera den nya regeringen , men här yppas inte ett ord om de bakomliggande orsakerna till fascismens uppgång .
denna framgång kan förklaras av förvirringen bland de folk som fallit offer för penningdyrkan och av de ledande klassernas val att främja en kraftig åtstramning , för att hela tiden kunna driva svångrems- och avregleringspolitiken ett steg längre .
för att opponera oss mot det främlingsfientliga talet hos en diktatorlärling som längtar tillbaka till det tredje riket , är alla tillfällen bra för att uttrycka vår solidaritet med de antifascistiska österrikarna .
därför kommer vi att rösta för denna resolution , trots de hycklande hänvisningarna till en &quot; europeisk demokratisk modell &quot; , som mer påminner om en fästning där man jagar , utvisar och låser in dem som lever under illegala förhållanden , när man inte sätter dit tonåringar .
- ( de ) jag har just röstat mot resolutionsförslaget om österrikes situation i betraktande av en möjlig regeringsbildning mellan österrikiska folkpartiet ( övp ) och österrikiska liberala partiet ( fpö ) .
jag håller det för kontraproduktivt att höja jörg haiders anseende som &quot; europas syndabock &quot; - en allvarlig nynazist och ledande rasist .
givetvis instämmer jag på intet sätt i denne högerpopulists publicerade uttalanden och fördömer på det starkaste all främlingsfientlighet och varje ansats till bagatellisering av hitler-regimen .
jag befarar dock att en blott och bart emotionellt präglad reaktion från europa på vad som sker i österrike kommer att mångfaldiga haiders anhängare .
europeiska unionen får inte skänka honom en pr-effekt som annars inte kan fås för pengar .
fpö : s styrka kan härledas till svagheten hos dem som hittills har regerat . här bär de österrikiska socialisterna huvudansvaret .
först efter att utan framgång ha propagerat hos fpö för accepterandet av en minoritetsregering och uppenbarligen förgäves ha erbjudit fpö ministerposter påbörjade österrikiska socialdemokratiska partiet ( spö ) sin massivt förda kampanj mot haider .
den hotande maktförlusten döpte de om till en &quot; heroisk kamp för upprätthållandet av värderingar &quot; och helt enkelt ett omedelbart förestående &quot; avgörande mellan demokratins vara eller icke vara &quot; .
detta är en smädelse mot väljarna i mitt grannland , vilken jag inte kan ställa upp på .
vi tyska kristdemokrater valde en annan strategi i kampen mot extremister och tog i klartext avstånd från dem .
vi avslöjade de innehållsliga bristerna hos rep ( &quot; die republikaner &quot; ) , vilka visade sig vara nationalistiska , främlings- och minoritetsfientliga .
i dag saknar rep representation i de flesta kommunalparlament .
den tyska vägen är ingen garanti för att denna radikala rörelse inte växer sig stark på nytt .
den kan inte tillämpas var som helst , eftersom varje medlemsstat har sina egna villkor .
övp ( österrikiska folkpartiet ) , som man inte längre kan ignorera ens på europeisk nivå , vågar sig på försöket med en koalition , för det österrikiska styrets skull .
detta kan lyckas endast om man träffar överenskommelser som på ett övertygande sätt bottnar i viljan att upprätthålla demokratiska grundläggande värderingar .
rådet har blandat sig i oöverlagt , utan att invänta resultaten av koalitionsförhandlingarna eller ett regeringsprogram .
detta fördömande är precis lika litet acceptabelt som hotet om att bryta kontakterna med republiken österrike
en väl befäst demokrati kräver att man är vaksam och inte blundar med ena ögat .
vi måste reagera offensivt och med argument mot radikala personer såväl från höger som från vänster .
jag skulle ha önskat mig samma häftiga europeiska protest när socialisterna såg sig redo att göra gemensam sak med efterföljarna till den människoföraktande och människoförföljande regimen i ddr .
sedan dess bildar de regering i olika tyska förbundsländer .
jag instämmer helt och fullt i de redogörelser som europeiska kommissionens ordförande prodi lämnade under dagens sammanträde .
han talade om vår plikt att inte isolera medlemsstater utan att göra allt för att knyta dem till gemensamma europeiska värderingar .
. ( fr ) jag har röstat emot den gemensamma resolutionen om situationen i österrike .
österrike är en fri , oberoende och suverän nation .
följaktligen kan varken rådet , kommissionen eller europaparlamentet blanda sig i en medlemsstats interna organisation .
valen i österrike har genomförts på ett fritt , regelmässigt och demokratiskt sätt .
därför är eu-institutionernas inblandning i det här landet oacceptabelt ; det är en kränkning av det europeiska fördraget ( artikel 7 i amsterdamfördraget ) .
likväl har dessa institutioner inte tvekat om att godkänna turkiets anslutning till europeiska unionen , samtidigt som man känner till att det förekommer kränkningar av de mänskliga rättigheterna .
ingen händelse av ett sådant slag har inträffat i österrike .
detta prejudikat , som skapats på initiativ av det portugisiska ordförandeskapet , är oroväckande för europeiska unionens framtid : dels avslöjar den politiska bannlysningen av österrike att likriktningen har ett oroande övertag , och dels kommer själva demokratins princip att förstöras om regeringarna i europeiska unionens medlemsstater i framtiden först måste - inte få folkets förtroende - utan nomineras av överstatliga organ .
kommer det att ens vara lönt att anordna val under sådana omständigheter ?
det är inte så man skapar förutsättningarna för att europas nationer skall kunna leva i harmoni och samarbeta för en gemensam framtid .
. ( fr ) den omröstning som just har ägt rum här är historisk , för det är första gången som vi med en så stor oro diskuterar den interna politiska situationen i en av våra medlemsstater .
jag tror det är lämpligt att frågan om institutionella principer och regler ställs åt sidan .
jag uppmuntrar rådet och dess ordförandeskap att fortsätta försvara unionens grundläggande värderingar .
och jag uppmanar kommissionen att vara mindre försiktig .
med denna resolution tar parlamentet sitt ansvar .
men samtidigt är den resolution som i dag antagits i mina ögon ett minimum minimorum , det minsta vi kan göra .
personligen har jag försvarat en ännu hårdare ståndpunkt och därmed stött ändringsförslagen 1 , 4 , 6 , 7 , och 8 , såväl som det muntliga ändringsförslag vilket föreslogs av socialistgruppen .
jag tror faktiskt att det är en nödvändighet att rådet endast accepterar tekniska förbindelser med företrädare för den österrikiska regeringen , där fpö-medlemmar kommer att ingå .
att låta jörg haiders parti ingå i en regeringskoalition kommer att banalisera extremhögern i europa , och utgör ett ytterst allvarligt prejudikat som skulle kunna dra med sig andra unionsmedlemmar eller kandidatländer .
här tar det österrikiska konservativa partiet ett historiskt ansvar .
det är våra grundläggande värden som står på spel ; i egenskap av européernas demokratiskt valda företrädare har vi inget val .
vi måste , våra väljare kräver det , vägra det oacceptabla .
när barbariets spöke dyker upp igen skall vi veta följande : &quot; att inte opponera sig är att kapitulera &quot; .
. ( fi ) jag röstade blankt vid omröstningen om resolutionen .
jag fördömer jörg haiders rasistiska och främlingsfientliga linje .
jag kan emellertid inte acceptera att eu : s organ gör en politisk intervention i en medlemsstats inrikespolitik .
därför kan jag varken godkänna punkt 4 i den gemensamma resolutionen eller rösta för resolutionen , inte ens mot extremhögern .
. det är uppenbart att de politiska ledarna i europa har rätt och skyldighet att reagera mot haider och hans parti .
de politiska ledarna i europa har rätt att uttala sin uppfattning om den politiska utvecklingen i ett annat medlemsland , på samma sätt som en statsminister kan uttala sig om rasistiska politiker i en kommun .
den finländska erfarenheten är emellertid att integrering är ett bättre sätt att bekämpa antidemokratiska krafter än att isolera .
därför röstade jag emot punkt 2 i resolutionen . detta förutsätter dock att alla parter respekterar mänskliga rättigheter .
eu-ordförandeskapets &quot; gemensamma reaktion &quot; på regeringsbildningen i österrike är juridiskt felaktig .
de 14 medlemsländernas reaktion saknar stöd i fördragen .
vi skall inte heller isolera de krafter i österrike som vill arbeta för mänskliga rättigheter .
trots dessa mina invändningar mot rådets agerande och min åsikt att det är bättre att verka för integrering än genom isolering , var det viktigt att visa klart var europaparlamentet står i frågor om rasism , varför jag röstade för resolutionen i slutomröstningen .
härmed avslutas omröstningarna .
jag förklarar europaparlamentets session återupptagen efter avbrottet torsdagen den 3 februari 2000 .
protokollet från sammanträdet torsdagen den 3 februari har delats ut .
jag förstår av er reaktion att många av parlamentsledamöterna inte fått protokollet , och det är självklart att ni inte kan justera ett protokoll som ni inte har fått .
jag föreslår därför att vi justerar det i morgon förmiddag , eftersom ni uppenbarligen inte fått det och det ber jag om ursäkt för .
justeringen av protokollet skjuts alltså upp .
fru talman ! rörande en ordningsfråga .
i förmiddags rapporterade bbc att en brittisk ledamot av europaparlamentet , som innehar en hög position inom sin delegation , fortsätter att erbjuda strategisk rådgivning till privata klienter , men inte meddelar i intresseregistret vilka dessa klienter är .
europas medborgare har rätt att förvänta sig att deras företrädare håller isär sitt privata vinstintresse från det allmännas bästa , men de kan bara vara säkra på att detta görs i varje enskilt fall om informationen både är tillgänglig för allmänheten och lätt åtkomlig .
fru talman ! eftersom dessa frågor för närvarande diskuteras i kvestorskollegiet , får jag be er att använda ert inflytande både för att se till att intresseregistret uppdateras och ändras för att omfatta fall av denna typ och , framför allt , för att se till att registret inte bara är tillgängligt för inspektion av denna kammare , utan att det också offentliggörs på internet ?
tack , herr davies .
jag skall titta på frågan med kvestorerna .
fru talman ! jag uttalar mig enligt artikel 9 i denna kammares arbetsordning och åsyftar samma fråga som togs upp av davies om de mycket allvarliga anklagelserna som uttalades på bbc i förmiddags .
jag skulle välkomna en försäkran från er att ni kommer att beställa en undersökning för att se till att de två ledamöter som nämndes i denna specifika bbc-intervju inte driver sina företag från detta parlament eller från parlamentets lokaler , eftersom detta i sanning skulle vara mycket allvarligt .
under årens lopp har de brittiska konservativas dubbelmoral gjort att det brittiska underhuset fått ett dåligt rykte , och det finns en verklig fara att ett sådant uppförande skulle få liknande effekter för detta parlament .
tack , herr murphy .
som jag sade till davies skall jag redan i kväll titta på frågan tillsammans med kvestorerna .
jag har redan skrivit till er vid ett flertal tillfällen om hur ordningsfrågor tas upp i kammaren .
jag undrar vilken ordningsfråga davies tog upp .
varför nämnde han inte att en av hans egna liberala kolleger också bedriver rådgivningsverksamhet som håller på att undersökas av bbc ?
skall denna kammare låta sin föredragningslista bestämmas av plumpa rapporter om ett program som grundar sina nyhetsinslag på lögner , eller skall den utföra ett seriöst arbete och ta itu med de utmaningar som europa står inför ?
kära kolleger ! det är självklart att kvestorerna som skall granska frågan inte enbart kommer att förlita sig på information som hörts i radion .
de kommer att gå igenom detta mycket noggrant .
fru talman ! jag tror att jag gör mig till tolk för ett stort antal kolleger i de flesta politiska grupperna när jag säger att det budskap som kommissionens ordförande framförde för en vecka sedan till den nya österrikiska förbundskanslern skapade obehag .
var det verkligen nödvändigt att säga , jag citerar : &quot; mina varmaste lyckönskningar följer er &quot; , eller &quot; jag betvivlar inte att ni kommer att fortsätta era föregångares engagemang när det gäller frihet och demokrati samt respekt för de mänskliga rättigheterna och grundläggande friheterna &quot; , eller &quot; jag ser fram emot ett fruktbart och konstruktivt samarbete &quot; ?
fru talman ! jag skulle vilja att prodi i morgon berättar för oss vad han ville eller inte ville ge för betydelse åt sitt uttalande så att ingen , absolut ingen , kan utnyttja detta minst sagt bisarra och olyckliga budskap , även mot prodis vilja , för att bidra till att banalisera den farliga politiska process som äger rum i österrike .
tack , herr wurtz . kära kolleger !
jag ber er att inte inleda någon debatt , det handlade om ett förslag som rör förfaranden .
jag vill erinra er om , herr wurtz , att vi i morgon träffar prodi som kommer att uttala sig om kommissionens program .
ni har naturligtvis full frihet att i era inlägg efter uttalandet fråga ut honom , på samma sätt som prodi har fullständig frihet att svara er .
jag föreslår att vi definitivt klargör denna fråga då , om ni och prodi vill det .
fru talman ! jag är mycket ledsen över att jag återigen måste besvära er med en punkt som jag redan tagit upp här två gånger tidigare .
jag har redan talat om för er ett antal gånger att vi för de nederländska kollegernas räkning gärna skulle vilja ha en nederländsk tv-kanal .
det finns nu 28 kanaler här i parlamentet , därav två grekiska , en portugisisk , en finsk och en belgisk , men fortfarande ingen nederländsk , däremot sju engelska , sex tyska och sex franska .
redan i september fick jag löfte om att det skulle finnas en nederländsk kanal i januari .
det är nu februari , och det finns fortfarande ingen .
jag skulle därför återigen vilja be er att vidta åtgärder för detta .
jag undrar vilken medeltida byråkrati det är som förhindrar att en nederländsk kanal överförs via satellit .
fru plooij-van gorsel ! jag är också besviken , eftersom jag själv var övertygad om att frågan hade lösts för länge sedan .
jag har noterat era budskap i frågan och jag tror att banotti har ett svar till er .
jag skall därför , om ni tillåter , lämna ordet till banotti så att hon kan svara er i form av ett förslag som rör förfaranden .
fru talman ! som min kära vän elly vet , kommer jag att göra allt för att se till att hon och mina nederländska kolleger blir nöjda .
jag kan i egenskap av kvestor med ansvar för denna fråga försäkra er om att vi haft tekniska diskussioner om de olika kanalerna på tv och radio , och jag har redan börjat skicka brev till kolleger i detta ärende .
om det nu kan lugna henne , har inte irländarna heller fått sin kanal ännu .
det verkar finnas svårartade tekniska problem , men vi arbetar verkligen på det .
tack för att jag fick möjlighet att reda ut detta .
jag är inte säker på att våra nederländska kolleger känner sig lugnade , eftersom våra irländska kolleger inte heller kan få in någon inhemsk kanal .
jag tror att vi måste titta på vad som kan göras så att alla kolleger kan se sin kanal .
tack , fru banotti , och övriga kvestorer , för era ansträngningar i ärendet .
fru talman ! jag ville säga till herr wurtz att kommissionens doktrin inte är bresjnevs doktrin om begränsad suveränitet och att vi inte , till dess att motsatsen bevisats , befinner oss inom ramen för artikel 6 och 7 .
österrike har därför fullständig rättighet att bilda en regering och kommissionens ordförande har fullständig rättighet , och till och med skyldighet , att framföra sina lyckönskningar till österrike .
wurtz kanske borde erinra sig att det inte var så länge sedan som kolleger i hans parti , franska kommunistiska borgmästare , skickade ut bulldozrar mot invandrarförläggningar i frankrike .
a ) sammanträdet den 14 till 18 februari 2000 i strasbourg beträffande onsdagen :
talmannen .
med tanke på att rådet inte kan vara närvarande onsdag kväll har flera grupper - europeiska folkpartiet , europeiska socialdemokratiska partiet , de liberala , de gröna och den enade vänstern - begärt att vi i en gemensam diskussion skall behandla rådets uttalande om den cypriotiska frågan och broks betänkande om föranslutningsstrategin för cypern och malta och flytta fram dessa punkter , liksom swobodas betänkande i föredragningslistan .
det skulle alltså innebära att vi på onsdagen har rådets två uttalanden om sammanhållningen mellan unionens politik och utvecklingspolitiken och om fn : s session om &quot; mänskliga rättigheter &quot; , följt av den gemensamma diskussionen om cypern och sedan om betänkandena från swoboda , frassoni och knörr borràs , samt rapporten från corrie .
vem vill lägga fram denna begäran i dessa gruppers namn ?
då ingen begärt ordet låter jag alltså begäran gå till omröstning .
( parlamentet biföll begäran . ) beträffande torsdagen :
när det gäller aktuella och brådskande frågor av större vikt har jag mottagit flera önskemål om ändringar .
när det gäller mänskliga rättigheter har jag mottagit två önskemål om tillägg : ett från den liberala gruppen om en underpunkt med beteckningen &quot; kambodja &quot; och ett från gruppen de gröna om en underpunkt med beteckningen &quot; pinochet &quot; .
som ni vet kan punkten &quot; mänskliga rättigheter &quot; inte omfatta fler än fem frågor .
förteckningen i det slutgiltiga förslaget till föredragningslista omfattar nu fyra frågor och vi kan därför bara lägga till ytterligare en .
vem vill lägga fram begäran om en underpunkt om kambodja för den liberala gruppens räkning ?
för den liberala gruppen är det av stor vikt att en diskussion om situationen i kambodja äger rum , och att det sker just nu . inte bara på grund av brevet som förenta nationernas generalsekreterare , kofi annan , skrivit till kambodjas regering för att den någon gång skall vida åtgärder för en särskild tribunal i syfte att ställa röda khmerernas ledare till svars , utan också för att hun sens regim , som uppenbarligen inte är nöjd med mordförsöken på oppositionsledaren sam raninsy , nu har kommit på att man kanske kunde upphäva hans parlamentariska immunitet för att han helt enkelt skall kunna ställas inför rätta .
världssamfundet har krävt att de skyldiga skall ställas till svars för det som sker i kambodja .
när allt kommer omkring var det vi som godkände valet i kambodja , vilket måste betecknas som ett av de största fiaskona på området valobservation .
det var bara parlamentet som kom ur detta med ett visst anseende i behåll .
jag tror att vi från parlamentets sida måste ta vårt ansvar även den här gången och göra ett uttalande om situationen i kambodja .
underpunkten kambodja läggs alltså till under punkten &quot; mänskliga rättigheter &quot; , vilket gör att begäran om en underpunkt rörande pinochet inte kan bifallas .
jag har också mottagit önskemål om att lägga till nya punkter i den aktuella och brådskande debatten om frågor av större vikt .
det handlar alltså inte längre om att lägga till frågor under rubriken &quot; mänskliga rättigheter &quot; , utan att lägga till nya punkter .
jag har mottagit tre önskemål : en första begäran från den enade vänstern om att lägga till en punkt &quot; moratorium om dödsstraff i förenta staterna och fallet med betty beets &quot; , en andra begäran från den liberala gruppen om att lägga till en ny punkt med beteckningen &quot; pinochet &quot; , och en tredje begäran från gruppen de gröna om att lägga till en ny punkt &quot; katastrofer : donaus miljö &quot; .
med tanke på den tid vi förfogar över , och eftersom vi som ni vet har ett uttalande från kommissionen om omstrukturering av företag , och den nuvarande förteckningen omfattar två punkter , kan vi alltså lägga till ytterligare två .
jag skall först ta begäran från gruppen den enade vänstern .
( parlamentet avslog begäran . )
vi går nu vidare till begäran från den liberala gruppen .
finns det någon som vill uttala sig för den ?
fru talman ! det är påfallande att europaparlamentet hittills inte har tagit ställning i fråga om det eventuella frisläppandet av pinochet trots de internationella häktningsorder som redan utfärdats .
med tanke på att den belgiska regeringens överklagande gillades förra veckan och med tanke på att beslutet i huvudsak ännu inte är fattat är det viktigt att parlamentet äntligen ger en ordentlig signal , en signal som borde innehålla att ingen kan undkomma en rättvis rättegång .
det är otänkbart att europaparlamentet , som med rätta ägnar så mycket uppmärksamhet åt respekten för de mänskliga rättigheterna , inte skulle göra något tydligt uttalande i detta fall .
fru talman ! detta är en fråga som är alldeles för allvarlig för att i nuläget behandlas som ett brådskande ärende .
för det första har europaparlamentet redan uttalat sig om general pinochet , men förutom det måste vi nu påminna oss vissa saker .
den första är att detta är ett ärende som är sub iudice i flera europeiska länder , och jag påminner kollegerna om att det ännu inte existerar ett europeiskt straffrättsligt område och inte heller ett europeiskt rättsområde .
vi är för den internationella brottmålsdomstolen , men den finns inte ännu .
för det andra finns det för närvarande en demokratiskt vald regering i chile , under ledning av ricardo núñez , vars första uttalande varit att alla som begått brott av detta slag skall ställas inför rätta . och jag påminner mig att den chilenska rättvisan , som är oberoende , för närvarande går igenom 60 stämningsansökningar mot general pinochet och hans brott mot mänskligheten .
jag anser att frågan är så viktig att vi bör följa den , men inte att vi skall lösa den med hjälp av förfarandet för brådskande ärenden .
vi är för att rättvisa skipas i denna frågan , men vi tror inte att det här är det lämpligaste sättet .
( parlamentet avslog begäran . ) talmannen .
vi kommer nu till den tredje begäran som är &quot; miljökatastroferna i donaus vatten &quot; , en begäran från gruppen de gröna .
finns det någon ledamot som vill lägga fram denna begäran ?
fru talman ! jag vill bara be kammaren att stödja detta förslag , eftersom det har varit väldigt många omflyttningar i denna föredragningslista .
det är ett ganska kort ärende , men det är extremt viktigt att det passerar parlamentet nu , och att det inte blir några förseningar .
det handlar nämligen om förfalskningar av euron , vilket är ett ärende som är väldigt brådskande .
vi har försökt driva igenom detta .
jag vore därför väldigt tacksam om kammaren skulle kunna stödja detta förslag .
beträffande fredagen : talmannen .
när det gäller fredagen har vi på förmiddagen en muntlig fråga om posttjänster och europeiska socialdemokratiska partiets grupp begär att resolutionsförslagen skall gå till omröstning direkt efter debatten och inte i bryssel , såsom föreslagits i det slutgiltiga förslaget till föredragningslista .
vill någon kollega yttra sig för pse-gruppen och lägga fram denna begäran ?
fru talman ! jag ber min vän enrique barón om ursäkt , men jag skulle vilja uttala mig emot detta förslag .
jag är till och med förvånad över att det dyker upp , eftersom vi hade kommit överens om detta efter diskussion i talmanskonferensen .
fru talman ! jag tror att ert förslag att dela upp det hela med debatt på fredag och omröstning senare är klokt .
skälet är följande : frågan berör inte mindre än 1 800 000 löntagare inom europeiska unionen .
vi har ett direktiv .
det är inte gammalt , det härrör från 1997 .
att inför ett nytt direktiv besluta om den framtida inriktningen i all hast , utan att ha tid att rådfråga fackföreningarna eller diskutera med samtliga parter på arbetsmarknaden , tycker jag strider mot den anda som vi vill ingjuta i debatten om frågor som direkt berör arbetsmarknadens parter .
jag är alltså för att vi behåller den ursprungliga uppdelningen : debatt på fredag , omröstning senare .
fru talman ! det är tydligen så att jag är skyldig wurtz en förklaring , och jag skall ge hela parlamentet den .
vi hade nått denna principöverenskommelse i talmanskonferensen .
jag visste inte då att kommissionär bolkestein skulle komma nästa vecka för att tala om denna fråga i utskottet för regionalpolitik , transport , och turism .
i min grupp har vi diskuterat frågan och , med beaktande av det nuvarande läget för hela integrationsprocessen av marknaden och avregleringen av en så känslig fråga , anser vi att det är lämpligt att parlamentet gör ett första uttalande , oberoende av vad det gör i framtiden , så att kommissionär bolkestein kan notera detta och för att ge en inriktning till debatten nästa vecka .
fru talman ! jag vill helt enkelt be kollegan wurtz att läsa igenom vad det här handlar om .
det är inte fråga om någon innehållslig kontrovers utan endast om frågesatsen : när skall kommissionen , efter att nu ha haft ett och ett halvt år på sig , äntligen vara i stånd att lägga fram direktivet ?
vad vi vill med resolutionen är bara att de utsatta tiderna skall hållas , och då är det viktigt att vi agerar så snabbt som möjligt .
därför vill jag stödja socialdemokraternas förslag att genomföra omröstningen på fredag .
fru talman ! cederschiöldbetänkandet avfördes ju från torsdagens föredragningslista .
därmed torde vi få litet tid över på torsdag .
eftersom vi , med hänsyn till det stora antal frågor som skall avhandlas på en och en halv timme , ju har mycket knappt om tid för de brådskande ärendena vill jag bara fråga sessionstjänsten om man inte kan undersöka huruvida vi kan få en halvtimme extra för de brådskande ärendena för att få talartiden att räcka .
det förefaller mig över huvud taget som om fördelningen av sessionstiden de senaste veckorna har varit mycket kaotisk .
det rådde stor tidspress under talartiderna , men så plötsligt hade vi en till en och en halv timme över förra torsdagen , då inget ämne fanns upptaget på föredragningslistan och vi blev tvungna att vänta på omröstningen .
på fredag i denna vecka har vi ett en fråga .
det är faktiskt absurt .
jag vill verkligen be om en granskning av hur ekonomiskt sessionerna planeras .
det är fullständigt möjligt : låt oss därför se om vi kan förlänga tiden för de brådskande frågorna med en halvtimme , eftersom cederschiölds betänkande utgår .
det är vad det handlar om , och enbart detta .
fru talman ! jag skulle vilja göra ett inlägg om en punkt på föredragningslistan för onsdagen , som ni inte tagit upp .
jag förstår att det inte är en polemisk fråga att uttalandet om 50-årsdagen av genèvekonventionerna inte innefattas i rådets uttalande om nästa möte i förenta nationernas kommitté för mänskliga rättigheter och att detta uttalande , för att utformas på ett ädelt och högtidligt sätt överlämnats till plenum i mars .
jag förstår att det finns en överenskommelse om detta .
fru talman ! under denna eftermiddag i denna kammare har det hänvisats till en rad rapporter på bbc : s program today denna förmiddag , i vilket man hävdade att vissa av mina kolleger drev personliga lobbyföretag eller på något sätt missbrukade sin ställning som ledamöter av denna kammare .
detta är allvarliga anklagelser .
de är fullständigt osanna , ondskefulla , politiskt färgade och de uttalades trots vetskapen om att de var osanna .
vi skall vidta rättsliga åtgärder .
mina kollegers intresseregister är fullständiga .
om vi får vetskap om att någon ledamot av denna kammare eller dennes medarbetare samarbetat med bbc i denna röra kommer vi att avslöja dem , vilket drar skam över denna kammare .
det stämmer , vi är helt överens .
b ) sammanträdena den 1 och 2 mars 2000 i bryssel
hållbar stadsutveckling - landsbygdens utveckling - equal-initiativet
( fr ) fru talman , kära kolleger , herrar kommissionärer och ledamöter av utskottet för regionalpolitik , transport och turism ! jag har fått i uppdrag att upprätta europaparlamentets betänkande om programmet för gemenskapsinitiativet interreg iii .
när frågan överlämnades till utskottet granskade vi över 100 ändringsförslag och hittills har 17 ändringsförslag på nytt lämnats in , vissa av dem har redan lagts fram för kommissionen .
innan vi diskuterar innehållet i den resolution som jag lägger fram skulle jag vilja tala om vilka beståndsdelar jag beaktat och använt som riktlinjer för mitt arbete som föredragande .
till att börja med vill jag erinra om den roll som gemenskapsinitiativet interreg har , som grundades på principen om gränsöverskridande och innovation .
programmet är en drivkraft när det gäller utveckling och den europeiska dimensionen .
interreg är ett av de fyra gemenskapsinitiativ som planeras för perioden 2000-2006 och kommer att förfoga över det största totalanslaget , nämligen 4,875 miljarder euro , jämfört med 3,604 miljarder för närvarande .
initiativet interreg inrättades 1990 och bygger på strävan att förbereda de europeiska regionerna för ett europa utan gränser , inom ramen för den stora inre marknadens genomförande .
vid reformen av strukturformerna 1994 och 1996 införlivades nya områden i gemenskapsprogrammet interreg , vilka bidrog till att utveckla transeuropeiska nät för transport och energidistribution .
dessa program har främjat gränsöverskridande samarbete , liksom samarbete mellan länder och regioner inom europeiska unionen , genom att främja en balanserad utveckling av gemenskapsområdet .
programmet interreg iii är en fortsättning av detta arbete och europeiska kommissionen överlämnar i dag riktlinjerna för detta till oss , i enlighet med bestämmelserna i rådets förordning ( eg ) nr 1260 från 1999 om allmänna bestämmelser för strukturfonderna .
programmet är uppdelat i tre områden : område a gäller det gränsöverskridande samarbetet mellan territoriella myndigheter och gränsregioner inom och utanför europeiska unionen , utifrån gemensamma utvecklingsstrategier och där genomförandet faller under medlemsstaterna och de lokala och regionala myndigheterna , område b gäller samarbete mellan länder och mellan nationella , regionala och lokala myndigheter i flera medlemsstater eller kandidatländer , inom områden som fysisk planering , transport- och miljönätverk .
genomförandet av detta område är medlemsstaternas och de nationella myndigheternas ansvar , och område c , slutligen , som gäller samarbetet mellan olika regioner i medlemsstaterna eller tredje land , med hjälp av erfarenheter från område a och b , samt samarbete inom forskning och teknisk utveckling , ett ämne som skall fastställas tillsammans med europeiska kommissionen , som ansvarar för genomförandet .
det nya interreg-programmet beaktar man i den form det överlämnats till oss de behov som uppstår genom utvidgningen till länderna i central- och östeuropa och till öregionerna och de yttersta randområdena .
kommissionen föreslår att vi skall fördela interregs resurser enligt följande : mellan 50 och 80 procent till område a , 6 procent till område c och skillnaden , dvs. mellan 14 och 44 procent , till område b.
europeiska kommissionen fastställer förteckningen över stödberättigade regioner inom område a och b och stöder sig huvudsakligen på kartan över stödberättigade regioner under föregående programplaneringsperiod .
de yttersta randområdena kan åtnjuta stöd inom område b. kommissionen upprättar en ofullständig förteckning över prioriterade områden och stödberättigade åtgärder för område a , men en fullständig förteckning när det gäller område b. kommissionen förbehåller sig rätten att senare föreslå frågor som den anser viktiga för utbyte av erfarenheter och förstärkt samarbete mellan regioner inom område c.
förfarandet för att anta programmen fastställs genom den allmänna förordningen om strukturfonderna .
förslagen upprättas av medlemsstaterna och överlämnas för godkännande till kommissionen , som kontrollerar att de överensstämmer med de allmänna riktlinjer som fastställts .
dessa förslag måste innehålla ett antal beståndsdelar , en överblick över gränsöverskridande eller transnationella strategier och prioriteringar , en beskrivning över de åtgärder som krävs för att de skall kunna genomföras och en vägledande finansieringsplan .
jag hör till den stora majoritet av parlamentsledamöter som röstat för att programmet för gemenskapsinitiativet interreg skall bibehållas .
jag beklagar att parlamentet inte informerats om utvärderingen av det tidigare programmet - vilket skulle ha gjort det möjligt att göra de nya åtgärderna optimalt effektiva , men jag vet hur svår denna åtgärd är - jag beklagar också att tidsplanen varit extremt kort , eftersom texten granskades i utskottet den 24 november och 26 januari , och jag beklagar också att vare sig de representativa regionerna eller regionala organisationerna fått möjlighet att delta i utarbetandet av programmet .
genom att främja ett gränsöverskridande samarbete mellan länder eller regioner är detta tvärgående instrument själva inkarnationen av en europeisk regionalpolitik som främjar en harmonisk och balanserad politik för fysisk planering inom gemenskapen .
( de ) fru talman , ärade kolleger ! mitt equal-betänkande har karaktären av ett yttrande inom ramen för rådfrågningsprocessen för ett nytt gemenskapsinitiativ , vars mål det är att få till stånd ett transnationellt samarbete för att främja nya metoder för bekämpandet av diskriminering och ojämlikheter av alla slag på arbetsmarknaden .
betänkandet blev mycket kostsamt eftersom det även inbegriper yttranden från fyra andra utskott - från utskottet för industrifrågor , utrikeshandel , forskning och energi , utskottet för regionalpolitik , transport och turism , utskottet för kvinnors rättigheter och jämställdhetsfrågor samt utskottet för rättsliga frågor och den inre marknaden .
detta gemenskapsinitiativ är en efterföljare till de två föregångarna adapt och employment och förfogar över en betydligt mindre budget , nämligen runt 2,8 miljarder euro .
initiativet slår in på en helt ny väg , nämligen för att ta fram innovativa sysselsättningsmodeller för transnationella utvecklingspartnerskap på geografisk eller sektoriell nivå .
avsikten är tydlig : det skall utvecklas riktade projekt på transnationell nivå , projekt som orienterar sig efter de sysselsättningspolitiska riktlinjerna , dvs. sysselsättningsförmåga , företagaranda , anpassningsförmåga samt lika möjligheter för alla .
denna målsättning skall verkligen välkomnas , och den finner gehör även i kammaren .
equal skall härutöver mynna ut i de nationella sysselsättningsprogrammen samt genom dessa åtgärdsprogram möjliggöra kontroll av införlivandet .
detta är ett viktigt gemenskapsinitiativ , som tillsammans med de tre andra initiativen urban , leader och interreg finansieras genom strukturfonderna .
jag har i rapporten försökt reducera de våldsamma förvaltningskostnaderna samt utforma starten på partnerskapet för utveckling något mer öppet och flexibelt .
jag anser att det tekniska stödet är nödvändigt , men på grund av problemen med de tidigare byråerna för utbyte av information om tekniskt bistånd skall det inte bli något nybildande av dessa byråer innan parlamentets resolution föreligger , och därmed skall förhindras att det politiska ansvaret läggs över på tekniskt bistånd .
men icke desto mindre är det tekniska biståndet nödvändigt .
särskild uppmärksamhet skall även riktas mot spridningen av resultaten och mot det ömsesidiga lärandet genom best practice och mainstreaming .
det har varit min strävan att kunna garantera att betänkandet får ett så brett stöd som möjligt .
detta har gjort att antalet ändringsförslag har minskats - från över 100 i utskottet till 22 för plenum - och det har sålunda även blivit möjligt att finna talrika kompromisser .
i frågan om asylsökande har det likaledes gjorts en kompromiss .
för att vi även skall kunna utforma detaljerna här ber jag dock , fru talman , att omröstningen om equal-betänkandet genomförs först på onsdag i stället för i morgon .
det är viktigt för mig att gemenskapsinitiativet kan köras igång i tid , att betänkandet får ett övertygande stöd så att kommissionen också manas att ta hänsyn till europaparlamentets konstruktiva förslag , för anslagen till equal har hållits tillbaka av europaparlamentet just för att ledamöternas invändningar skall komma till uttryck i detta gemenskapsinitiativ .
därför är det också befogat att parlamentet insisterar på att ämnesprioriteringarna skall kunna ändras först efter att parlamentet har hörts på nytt .
equal skall , och det är min bestämda avsikt , göra rättvisa åt sitt namn .
genom det skall alla eftersatta grupper i europeiska unionen erbjuda samma chanser .
det skall förhindra att samhället faller isär .
det skall hindra utslagningen från att vara en del av vardagen .
alla skall erbjudas möjligheten att dra fördel av ett gemensamt initiativ , oavsett hur gamla eller av vilket kön de är och varifrån de kommer .
detta är min avsikt , och jag ber om ett övertygande stöd för betänkandet i kammaren !
fru talman ! det är i sig självt en prestation att vi har denna debatt om gemenskapens nya stadsmiljöinitiativ inom urban-programmet , och det är en prestation att jag är här i kväll , eftersom air france ställde in mitt flyg som skulle gå kl. 14.10 - men jag är här !
för bara ett år sedan när kommissionen utarbetade sina förslag kring agenda 2000 skar man ned stadsmiljöinitiativet .
ändå visste vi i egenskap av politiker att det fanns en underström av stöd för en fortsättning av detta initiativ under år 2000 .
parlamentet kan därför ta åt sig äran för att ha genomfört en framgångsrik påtryckningskampanj för att få tillbaka urban-programmet på dagordningen och få kommissionen och rådet att göra en kovändning .
stadsmiljöpolitiken har alltid varit högt prioriterad inom eu : s politik .
i min medlemsstat , t.ex. , håller vi på att utveckla ett strategiskt förhållningssätt genom en vitbok och en statlig stadsmiljögrupp håller på att undersöka de problem som finns i stadsmiljön .
i ett läge där 80 procent av befolkningen i europa bor i stadsområden , är det rätt och riktigt att vi hjälper våra mest eftersatta samhällen att ta itu med de alltför bekanta problemen med förfall , social utslagning , arbetslöshet , kriminalitet , drogberoende och alla de problem som har samband med detta .
i min hemregion , t.ex. , i manchester , har stadsmiljöinitiativet inom urban-programmet blivit en enorm framgång .
medel från programmet har investerats i ett av de mest förfallna stadsområdena i förenade kungariket , moss side .
&quot; the millennium youth park &quot; projektet hjälper till med att få unga personer intresserade av att rusta upp sitt eget grannskap och förutom stöd till mindre företag och socialpolitik , börjar vi se en återhämtning inom detta mycket eftersatta stadsområde .
arbetet med denna urban-dagordning togs sedan till andra delar av samhället med en aktiv kommunikations- och offentlighetskampanj på lokala stormarknader och berömda brittiska pubar .
det är denna typ av bra åtgärder som vi också vill skall utvidgas till hela eu när det rör kommunikation och offentlighet .
vad gäller de särskilda riktlinjer som styr initiativet , är de flexibelt definierade för att ge utrymme för lokal och regional mångfald .
vi håller med om att de bör vara vägledande till sin natur och låta en maximal flexibilitet se till att vi uppnår specifika programmål .
i utskottet förespråkar vi inte en minskning av antalet till 50 .
vi förespråkar en allmän minskning , men vi anser inte att den godtyckliga siffran 50 är den viktigaste faktorn .
vi borde i stället satsa på högkvalitativa projekt som kan fungera som en katalysator för förändring och förnyelse , som kan dra till sig investeringar rörande lån och riskkapital och åstadkomma en multiplikatoreffekt .
medlemsstaterna bör därför kunna föreslå ett skäligt antal områden inom det finansiella taket för sina anslag .
vid angivandet av lokala urban-program , måste vi verkligen ta hänsyn till lokala indikatorer och lokal statistik om eftersatthet och hälsotillstånd för att vi skall kunna ta itu med de värst drabbade områdena på ett mer effektivt sätt .
i förenade kungariket är det lokala eftersatthetskriteriet ett mycket bra exempel på en allmänt använd standard och statistik till hjälp för att bestämma inte bara stödprogram inom eu , utan också nationella och regionala stödprogram .
detta måste börja användas som ett instrument och en resurs , som ett komplement till eu-kriterierna .
jag vill be er att ta hänsyn till lokala indikatorer för att hjälpa oss med detta .
våra mest eftersatta stadsområden står inför en överväldigande mängd problem : hög arbetslöshet och ofta mycket dåligt betalda och osäkra jobb , fattigdom och social utslagning .
dessa problem förvärras ofta genom dåligt hälsotillstånd , dåliga bostäder och en kultur där drogberoende ingår .
det är därför vi har fått instabila samhällen som genomsyras av kriminalitet , narkotikahandel och gäng .
detta är alltför välbekant i många av våra stadsområden .
alla dessa komplexa problem undergräver livskvaliteten för de stadsboende , fast möjligheten finns i dessa områden att skapa tillväxt och välstånd .
detta är återigen skälet till varför jag i mitt betänkande har poängterat att åtgärder i samband med urban-programmet inte bara bör tillhandahålla en helhetslösning till ett enda problem : dessa områden lider inte av enstaka problem .
samhällena i stadsområdena bör i stället uppmuntras till att lägga fram integrerade handlingsplaner som kan hjälpa till med att lösa deras specifika stadsrelaterade problem , genom att använda eu-resurser som ett komplement till lokala åtgärder .
jag skulle vilja se att dessa åtgärder utökades till att omfatta hälsofrågor och åtgärder mot diskriminering , som fastställts i amsterdamfördraget .
gemenskapsinitiativet innebär gemenskapsengagemang .
några av de mest aktiva och engagerade krafterna för förändring inom våra stadsområden är de personer som bor där .
vi måste uppmuntra dem att delta i utformningen och slutförandet av projekt inom dessa program .
den tidtabell som föreslagits av kommissionen är därför mycket ambitiös .
det är bättre att ha kvalitetsprojekt med ett aktivt deltagande av gemenskapsgrupper , än att ha projekt som slutförs enligt tidtabell men utan lokalt deltagande .
kommissionen måste naturligtvis se till att det råder fullständig öppenhet rörande de urvalskriterier som används för de nya programinitiativen , men den måste också redovisa vilka rådgivningsnätverk som används för utbytet av bästa metoder .
detta är viktigt när det rör öppenhet och nätverkens övergripande effektivitet .
låt mig till sist betona att vi behöver lokalt engagemang för att kunna ta itu med de problem som det postindustriella samhället står inför .
vi måste använda oss av de arbetslösas inneboende kraft , ungdomarnas för litet använda färdigheter och de äldres erfarenheter för att kunna lösa dessa problem .
vi skall då kunna ersätta fattigdom , beroende och främlingsskap med rättvisa , initiativkraft och deltagande .
detta kommer att hjälpa oss att återställa eu : s trovärdighet och medborgarnas tro på att europeiska unionen kan få till stånd lokala åtgärder för att lösa lokala problem .
( it ) herr talman ! som föredragande mccarthy redan har påmint om kan urban verkligen betraktas som en seger för europaparlamentet som en följd av den debatt som pågick förra året om reformering av förordningarna .
som har sagts är syftet med urban att främja innovativa strategier till förmån för en ekonomisk och social nylansering av stadsområdena , också mot bakgrund av att 80 procent av europas befolkning är koncentrerad till städerna .
att skapa en positiv stadsmiljö ur socialpolitisk synvinkel innebär att förverkliga en politik som syftar till att skapa varaktiga arbetstillfällen , att bekämpa fattigdomen , att vidta åtgärder till förmån för låginkomsttagare , äldre och barn , etnisk och rasmässig integration , bättre möjligheter till delaktighet , en profilerad hälso- och sjukvårdspolitik som omfattar åtgärder för att förebygga drogberoende liksom en samordnad brottsförebyggande politik .
kommissionen tar i sitt meddelande hänsyn till behovet av angreppssätt som omfattar ett helt spektrum av ekonomiska och sociala infrastrukturåtgärder .
emellertid måste man komma ihåg att det förutom urban finns flera andra gemenskapsinstrument på det sociala området : innovativa åtgärder enligt europeiska socialfondens artikel 6 , pilotprojekt - framför allt den nya förberedande satsning på &quot; lokala sysselsättningsinitiativ &quot; , som europaparlamentet nyss införde i och med budgeten för 2000 - initiativen equal och interreg liksom mainstreaming av socialfonden .
som utskottet för sysselsättning och socialfrågor understryker i sitt yttrande måste alltså kommissionen ta hänsyn till synergieffekter i detta sammanhang och samtidigt undvika dubbleringar inom de finansierade projekten .
samtidigt som vi å ena sidan anser det nödvändigt att styrkommittéerna säkerställer att de olika insatserna är inbördes konsekventa och kompletterar varandra , uppmanar vi å den andra sidan kommissionen att öka informationsutbytet och samordningen mellan de avdelningar som berörs .
en sådan samordning är inte det enda som är viktigt , utan även utbytet och spridandet av erfarenheter och god praxis måste vara viktigt , vilket vi påpekar i vårt yttrande .
herr talman ! betydelsen av detta initiativ blir allt större allt eftersom de ekonomiska och sociala problemen förvärras i europas städer och allt eftersom invånarna i städerna känner sig allt med fjärmade från sina städers eller förorters förvaltning .
till denna situation kommer de sociala omstruktureringarna till följd av utvidgningen av europeiska unionen att komma till , och följaktligen måste vi i god tid ombesörja våra städers ekonomiska förnyelse och sociala sammanhållning .
dessa problem måste för övrigt bemötas även med tanke på städernas stora inflytande på de kringliggande regionerna , liksom även med tanke på deras historiska och kulturella roll .
för att våra ansträngningar skall lyckas , krävs det emellertid att alla medborgare engagerar sig och deltar samt att de mindre aktiva samhällsgrupperna och de grupper som drabbas särskilt hårt av den ekonomiska och sociala krisen aktiveras .
och här vill vi betona nödvändigheten av att kvinnorna , eller de aktörer som företräder kvinnorna , på ett balanserat sätt deltar i planeringen och genomförandet av urban-initiativets program .
vi i utskottet för kvinnors rättigheter och jämställdhetsfrågor betonar även nödvändigheten av att finansiera infrastrukturer som gör det lättare för kvinnorna att vara yrkesverksamma , huvudsakligen med avseende på en harmonisering av yrkes- och familjeansvaret , och bredare infrastrukturer som främjar generationernas solidaritet , den sociala solidariteten .
om detta initiativ genomfördes på ett effektivt sätt , skulle det kunna få en multiplikatoreffekt , eftersom det skulle kunna stimulera till liknande åtgärder på regional och lokal nivå . initiativets politiska betydelse skulle då bli ännu större , eftersom kvinnorna behöver känna påtagliga resultat av den europeiska politiken i sina vardagliga liv .
( de ) herr talman ! vi har i vårt utskott välkomnat det faktum att kommissionen har föreslagit att urban-programmet skall prioritera en bättre integrering av lokala gemenskaper och etniska minoriteter liksom höjningen av säkerheten och förebyggande åtgärder mot kriminalitet .
vi har i utskottet ansett det nödvändigt att ett ekonomiskt och socialt återupplivande av stadsområden åtföljs av en atmosfär med tolerans gentemot minoriteter , så att åtgärder avsedda att minska rasism och främlingsfientlighet blir ett integrerat inslag i de program som skall finansieras inom ramen för urban .
vi har ansett att en central uppgift när det gäller återupplivandet av stadsområden är att höja medborgarnas känsla av trygghet och därmed att bekämpa vardagskriminaliteten i städerna .
utskottet har konstaterat att en nytänkande och effektiv kriminalitetsbekämpning liksom förebyggandet av kriminalitet kräver åtgärder som differentieras på kommunal nivå - hit hör att förebyggandet av kriminalitet tas med i stadsplaneringen , åtgärder för att förebygga ungdomsbrottslighet , återanpassning av förbrytare liksom modeller för ett verkningsfullt samarbete mellan olika aktörer på lokal nivå , t.ex. polis , rättsväsende eller sociala instanser .
i utskottet har vi enhälligt ställt oss bakom rekommendationen , eftersom vi var mycket angelägna om att just urban - som i tidigare skeden har varit ett så framgångsrikt gemenskapsinitiativ - får en fortsättning , för vi utgår ifrån att vi endast med hjälp av dylika program inom europeiska unionen kommer att lyckas förverkliga en fredlig samexistens på sikt för alla invånare i europeiska unionen .
det är av den anledningen som vi varmt välkomnar denna typ av program .
ättning och socialfrågor . ( de ) för det mest omfattande av de fyra gemenskapsinitiativen , nämligen interreg iii , vill jag föra fram önskemålen från utskottet för sysselsättning och socialfrågor .
det måste finnas möjlighet att satsa stort även på sociala åtgärder när det gäller interreg iii .
med tanke på att 50 procent av arbetslösheten i unionen till väsentliga delar är strukturellt betingad och med tanke på den särskilt känsliga situationen i gränsområdena - jag pekar endast på möjliga oönskade migrationsrörelser - är detta inte bara förnuftigt , utan nödvändigt .
nu tycks också de stödåtgärder som anförs i bilaga ii till programinriktning a vara lovande i detta hänseende .
men i kommissionens meddelande saknas det faktiskt helt och hållet bestämmelser för medlemsstaterna som omfattar dessa integrerade satsningar på social- och sysselsättningspolitiska aspekter .
därför vill jag särskilt betona ett ökat insättande av yrkesutbildningsåtgärder , i synnerhet i områden med hög långtids- och ungdomsarbetslöshet .
inriktning b bör likaledes vara öppen för sysselsättningspolitiska stödåtgärder , speciellt i samband med strategin för att föra fram medlemskandidaterna .
när det gäller de sysselsättningspolitiska åtgärderna ser jag det rent generellt som en nödvändighet att den gemensamma samarbetskommittén tillsätts regionalt därför att närheten och den nödvändiga sakkunskapen som rör dessa åtgärder bara finns på regional nivå och därför att det skall förhindras att åtgärderna blir verkningslösa .
att förvaltningskostnaderna för interreg iii - som jag ser det - fortfarande är för höga kan vi alltid kritisera , det måste vi också hela tiden göra , även om jag nästan börjar tro att detta är oundvikligt i kommissionens stödprogram .
jag vill dock påpeka att det är ödesdigert just här .
just vad gäller sysselsättningspolitiken bör vi eftersträva så enkla åtgärder som möjligt för att den sociala dimensionen i europeiska unionen återigen skall ges den tyngd som den förtjänar .
utskottet för regionalpolitik , transport och turism tittade bl.a. på meddelandet om leader + och beslutade att stödja decentraliseringsprocessen i hanteringen av åtgärder . man ansåg att en sådan process kan vara effektiv om man uppfyller två villkor : att de lokala aktionsgrupperna är representativa för lokalsamhällets allmänna intressen och att kommissionens kontrollmekanismer används för att undvika att de territoriella och lokala myndigheterna använder medel från leader + för att bibehålla organisationer och civila grupper vinklade till myndigheten .
det begärs att man i de organ som fattar beslut om projekten garanterar en likvärdig representation av tre komponenter : de politiskt valda och offentliga myndigheter , företagen och de ekonomiska parterna , samt arbetsmarknadens parter , inklusive fackföreningar och frivilligorganisationer .
särskilt understryks att det skall vara en jämn könsfördelning i alla dessa organ .
man understryker dessutom att huvudsyftet är att främja strategier för en hållbar utveckling , vars positiva effekter skulle sträcka sig över ett bredare geografiskt område än själva lokalsamhället , och man anser det således vara lämpligt att projekten innefattas i utvecklingsprogrammen , inklusive mål 1 och 2 samt i planerna för den fysiska planeringen i de regioner och länder där de lokaliseras .
man gläds åt att leader + kan användas i alla landsbygdsområden i unionen , men man beaktar dock att det är nödvändigt med en koncentration av gemenskapsresurserna till de mest missgynnade regionerna för att underlätta den socioekonomiska sammanhållningsprocessen i unionen , utan att de statliga myndigheterna styr dessa medel mot syften som inte har med sammanhållningen att göra .
utskottet är av den uppfattningen att man för de projekt som finansieras inom ramen för åtgärd 1 borde värdera potentialen för en endogen utveckling , som i synnerhet stöds på lokala traditioner , tekniker och vanor , på specifika produktioner och på en hållbar energiutvinning .
utskottet stöder kommissionens förslag att koncentrera åtgärderna till ett reducerat antal valda områden och är av den uppfattningen att med hänsyn tagen till de olikheter som finns i många samhällen på landsbygden skall det demografiska minimitaket för att välja ett projekt minskas till 10.000 invånare .
man anser att det är nödvändigt att samordna utvecklingsmålen och mekanismerna för hantering av åtgärderna 2 och 3 som finansieras av leader med övriga åtgärder som finansieras med hjälp av andra gemenskapsprogram för samarbete och interregionala och internationella partnerskap , som interreg , sapar , phare , tacis och meda inom samma områden .
( de ) ärade herr talman , ärade fru föredragande , ärade kolleger ! innan jag närmare går in på equal-betänkandet vill jag säga något principiellt om de riktlinjer för sysselsättning som ligger till grund för betänkandet .
de grundläggande målen med en gemensam sysselsättningspolitik för eu har där fastställts till att gälla bland annat sysselsättningsförmåga , företagaranda och anpassningsförmåga .
dessa mål syftar uppenbarligen till att göra arbetstagarna så nyttiga och exploaterbara som möjligt för näringslivet .
ett försök att verkligen avveckla diskriminering på ett effektivt och långsiktigt sätt skulle emellertid behöva ha människors självbestämmande som mål .
först då handlar det inte längre endast om ekonomisk användbarhet , utan om ett jämlikt sätt för människor att gestalta sina liv .
likväl har stenzels betänkande utvecklats bra , åtminstone det som rör de fastställda riktlinjerna .
alla asylsökande och flyktingar skall uttryckligen omfattas av programmet , vilket emellertid borde vara en självklarhet .
ändå har de konservativa i utskottet röstat emot detta .
till dessa personer har jag en fråga : är målet med er politik att marginalisera människor ?
vad är det för idé som ligger bakom att förvägra människor arbete när de vill arbeta ?
står inte det i rak motsats till riktlinjen &quot; sysselsättningsförmåga &quot; ?
det är också värt att nämna att det här handlar om ett mainstreaming-program , för betänkandet är förenat med vissa brister .
sålunda betonas särskilt aspekten att kvinnor skall beredas bättre möjligheter på arbetsmarknaden genom att fler förskolor skall byggas .
den som låter männen klättra ostört uppför karriärstegen och enbart bekymrar sig om daghemsplatser utan att bekämpa den ojämna fördelningen av det reproduktiva arbetet , han och dessvärre även hon har inte förstått vad mainstraming är !
herr talman , ärade damer och herrar ! utskottet för regionalpolitik , transport och turism har vid de avslutande överläggningarna enhälligt , dock med en nedlagd röst , godkänt föreliggande yttrande om equal-betänkandet .
detta placerar jag medvetet först i min redogörelse för att tydliggöra att det faktiskt föreligger en motsättning mot det ansvariga utskottet för sysselsättning .
att samtliga grupper har godkänt yttrandet kan förklaras av de slutsatser som är ägnade att koppla samman regional- och transportpolitiska frågor liksom turismfrågor med bekämpningen av diskriminering och ojämlikheter av alla slag på arbetsmarknaden .
ledamöterna i utskottet för regional ser naturligtvis även en rad kritiska moment i kommissionens förslag , för det första har exempelvis den tematiska orienteringen för utvecklingspartnerskapens agerande inte fastställts i tillräcklig utsträckning ; för det andra återstår det fortfarande för kommissionen att utarbeta strikta urvalskriterier för utvärderingen av projektförslagen ; för det tredje befarar man för höga förvaltningstekniska kostnader för projektledningen via kommissionen liksom instanserna för det tekniska biståndet .
därför skall en övre gräns dras för förvaltningsuppgifterna .
utskottet har dragit slutsatser av dessa kritiska anmärkningar .
särskild vikt lägger vi vid kopplingen mellan skapandet av nya arbetstillfällen för socialt missgynnade och utslagna personer , inom turismen såväl som inom de små och medelstora företagen , och stödet för bildandet av små och medelstora företag med hänsyn till den nödvändiga ekonomiska strukturförändringen .
sammanflätningen av aktiviteterna inom gemenskapsinitiativen och de europeiska sysselsättningsinitiativen är ett grundläggande krav och en avgörande förutsättning för att equal-programmets olika uppgifter skall kunna fullgöras .
vi stöder eftertryckligen det innovativa försöket att bilda internationella utvecklingspartnerskap och att organisera utbytet av erfarenheter på europeisk nivå som en integrerad beståndsdel i equal-programmet .
den speciella målsättningen att nå europeisk framgång lyfter upp det regionala samarbetet till europeisk nivå samtidigt som samarbetet mellan de mest skilda regionala aktörer bibehålls .
detta är bra , och därför har vi också rekommenderat det .
herr talman , bästa föredragande , bästa åhörare ! jag tackar föredragandena som på kort tid åstadkommit sakkunniga betänkanden .
i min grupp har man dock kritiserat tidpunkten för utskottets förberedelsearbete .
betänkandena är försenade , dessutom drevs behandlingen åtminstone i utskottet för regionalpolitik , transport och turism med en stor brådska .
på så vis missade man ett bra tillfälle att debattera resultatet av tidigare program , god praxis och även brister .
vår grupp betonar i samband med interreg-programmet den gränsöverskridande verksamheten och i synnerhet det samarbete som sträcker sig utanför unionens gränser .
viktiga regioner är bland annat balkan och regionerna vid adriatiska havet , men enligt min mening bör man inte heller glömma samarbetet med ryssland .
vår grupp vill på nytt lyfta upp den praktiska kontrollen av fonderna och framhåller bland annat vikten av en bättre samordning mellan interreg- , tacis- , ispa- och phare-programmen .
i dag saknas denna samordning , och kommissionen har fortfarande inte lagt fram exakta förslag för att förbättra samordningen .
vi här i parlamentet förväntar oss att kommissionen så snabbt som möjligt skall lämna en noggrannare redogörelse av frågan inför vårt utskott .
när det gäller det praktiska genomförandet är det av avgörande betydelse att få med sig lokala företag , organisationer och andra aktörer .
erfarenheten har visat att det i samarbetsprojekten behövs bättre planering , noggrannare uppföljning och genomförande som leder till bättre resultat .
projekten har ofta stannat halvvägs och effektiviteten försvunnit i förvaltningen och byråkratin .
man måste också kräva av samarbetspartner att de förbinder sig till projekten och uppfyller sin egen del .
vår grupp lägger på nytt fram några ändringsförslag som avslogs vid utskottsbehandlingen .
jag tar här upp urban-betänkandet där föredraganden i motiveringar på ett förtjänstfullt sätt behandlat det minimibelopp på 500 euro per invånare som ingår i kommissionens riktlinjer .
det fungerar inte som ett mekaniskt mål utan det måste kunna anpassas efter förhållandena i målområdet .
detta är en så viktig synpunkt att det måste lyftas från motiveringar till slutsatser .
herr talman , kära kolleger ! interreg är en av de mest europeiska av alla strukturfonder .
här skall projekt stödjas inte bara i en region , i ett land , utan i angränsande regioner i två eller flera länder .
tyvärr gäller detta endast en del av pengarna , nämligen endast för gränserna inom eu .
men just de regioner som gränsar till tredje land är de som behöver ett fungerande verktyg för ett gränsöverskridande samarbete .
förordningen ger sken av att det också skulle förhålla sig så .
men så förhåller det sig inte . det förhåller sig nämligen så att kommissionen inte har ändrat förordningen på flera år , trots att parlamentet kräver detta sedan länge .
för regionerna innebär det i praktiken att det den närmaste tiden återigen degraderas till att likna västtysklands tidigare stödåtgärder till förfallna områden längs gränsen mot östtyskland .
parlamentet har sedan 1996 krävt att en gemenskapsfond bildas för samarbetet med tredje land för att lösa problemen .
ingenting har hänt !
man drar ytterligare ut på tiden med problemen , på berörda regioners bekostnad .
parlamentet kräver på nytt en förbättring och ett gränsöverskridande samarbete , och vi förväntar oss att en gemenskapsfond bildas och att förordningen ännu en gång ändras i samarbete med övriga kommissionärer .
vi vill ha ett medborgarnas europa och inte ett byråkraternas europa !
herr talman ! en tredjedel av europeiska unionens pengar stoppas in i fonder för allehanda utvecklingsändamål .
min grupp anser att det är utmärkt om detta leder till att man arbetar bort eftersatta regioner , städer eller befolkningsgrupper eller att hälsan och miljön förbättras .
det är en fråga om solidaritet och utveckling .
men att dela ut alltmer pengar är ingen garanti för att de också används på ett allt bättre sätt .
kommunerna och regionerna där pengarna hamnar har med tiden fått praktisk erfarenhet .
de konstaterar att det är ytterst svårt att använda pengarna till de ändamål där de allra bäst behövs .
det brukar för det mesta gå bra med allt som faller under ekonomisk tillväxt och infrastruktur , men det är ofta inte helt säkert att sociala ändamål och miljösyften blir godkända .
eftersom det råder stor osäkerhet om hur reglerna skall tolkas hyr kommuner och regioner nu in dyra byråer .
dessa sakkunniga får till uppgift att göra en uppskattning av i vilken grad europeiska kommissionens tjänstemän är beredda att godkänna planerna .
i vissa fall får jag intryck av att det inte handlar om solidaritet eller om att lösa de mest akuta problemen , utan om att upprätthålla befintliga intressen och om propaganda för europeiska unionens välsignelser .
det förefaller som om den viktigaste målsättningen på detta område har blivit att snickra ihop och måla propagandaskyltar där det står att ifrågavarande projekt medfinansieras av europeiska unionen .
det är för mycket pengar som går till spillo på propaganda och utredningsbyråer , på överläggningar och kontroll , och mycket pengar går tillbaka till det land som de kom ifrån .
efter den planerade anslutningen av nya medlemsstater med 100 miljoner invånare , där välfärdsnivån ligger på en tredjedel till två tredjedelar av genomsnittet för dagens medlemsstater i europeiska unionen , kommer detta slöseri att skapa ännu fler nackdelar .
i utskottet för regionalpolitik , transport och turism var gruppen enade vänstern överens med föredraganden av yttrandet om leader , nogueira román .
med rätta konstaterade denne att det inte ligger något positivt i att sprida alla dessa medel över alla landsbygdsområden .
i valet mellan innovationsprojekt och att koncentrera pengarna till att bekämpa eftersatthet väljer vi det sistnämnda eftersom detta ger det största bidraget till jämlikhet .
innovation i områden där det redan går bra ger ju redan avkastning och kommer att äga rum även utan europeiska bidrag .
ytterligare en punkt att uppmärksamma är risken för maktmissbruk och svågerpolitik inom regionala och kommunala förvaltningar .
tonvikten ligger på lokala grupper där myndigheter , organisationer och vinstinriktade företag samarbetar .
diskussionen har handlat om den fördelningsnyckel som skall tillämpas i sammanhanget .
här har bland annat en variant varit på tal som för tankarna till den nederländska &quot; poldermodellen &quot; , det strukturellt organiserade samarbetet mellan stat , fackförbund och företagarorganisationer .
låt oss inte glömma bort att val till kommunfullmäktige och regionala församlingar hålls för att företräda hela befolkningen .
egentligen borde det vara så att dessa organ gör en avvägning och då tar hänsyn till fackföreningsrörelsens och miljörörelsens önskemål .
min grupp motsätter sig inte att fackföreningsrörelsen och miljörörelsen , vars insatser i samhället vi anser vara viktiga , tilldelas en egen tydlig roll .
det kan förekomma att deras insatser förbigås på grund av lokala förvaltningar som fungerar kortsiktigt eller som inte fungerar tillräckligt demokratiskt .
men det faktum att vi nu måste vara rädda för maktmissbruk och svågerpolitik antyder att demokratin tyvärr ännu inte fungerar optimalt .
en invändning är att de valda organens begränsade roll medför att företag får mer inflytande .
så länge ekonomin inte vilar på demokratiska avvägningar av allas behov i stället för vinstintresset för några få är det tveksamt om demokratin fungerar bättre under inflytande från företagare än under inflytande från kommunfullmäktige .
för oss handlar det om &quot; en människa , en röst &quot; i stället för &quot; en aktie , en röst &quot; .
herr talman ! det finns ekonomiska gränser inom europeiska unionen och vid rådande tidpunkt fungerar den inre marknaden med fri rörlighet för varor , personer , tjänster och kapital helt och fullt .
men om den inre marknaden skall kunna fungera effektivt och om den gemensamma europeiska valutan skall bli framgångsrik , är det viktigt att alla regioner i europa - det finns över 100 - kan konkurrera ekonomiskt inom denna mycket utmanande miljö .
vissa områden i europeiska unionen är ekonomiskt sett mycket starka och överskrider mycket tydligt den genomsnittliga inkomsten per capita .
det finns fattiga regioner i unionen som måste få stöd från gemenskapen för att förbättra strukturerna hos sina ekonomier , så att de kan konkurrera inom europeiska unionens struktur .
om vi tittar på eu : s budgetplan mellan 1989 och 1993 , och 1994 och 1999 , är det därför vi kan konstatera att en så stor andel av eu : s budget avsattes för förvaltningen av europeiska regionala utvecklingsfonden och europeiska socialfonden .
det finns dubbla problem som fortfarande återstår för många europeiska regioner : för det första har vi bristen på lämplig infrastruktur vad gäller vägar , vattenreningsanläggningar och transportnät i detta sammanhang ; för det andra har vi behovet av att få igång initiativ för att bekämpa ungdoms- och långtidsarbetslöshet , som är ett ständigt socialt problem i många stads- och landsbygdsområden i europa .
det måste alltid finnas ett engagemang för att se till att vi inte bara bygger ett städernas europa .
vi måste se till att det sätts igång sysselsättningsskapande initiativ som främjar sysselsättningen inom sektorn för små och medelstora företag , även på den europeiska landsbygden .
de huvudsakliga aspekterna av debatten denna kväll har samband med funktionen hos gemenskapsinitiativen , dvs. de nya interreg iii- , equal- och leader + -initiativen .
mellan dessa tre program måste det finnas en tydlig demonstration av eu : s engagemang för främjande av en gränsöverskridande utveckling , kampen mot problemen i samband med långtidsarbetslöshet och stöd till program för landsbygdsutveckling .
herr talman ! det finns en hel del städer i europeiska unionen som har att kämpa med det underläge de befinner sig i .
det finns inte alltid tillräckligt med medel tillgängliga inom medlemsstaterna för att ta itu med detta på ett effektivt sätt .
därför är det meningsfullt att europeiska unionen fortsätter att stödja medlemsstaterna och , om så behövs , ger kompletterande stöd inom ramen för urban .
kommissionens förslag beträffande urban innehåller en nedskärning för de kommande sju åren , både i fråga om gemenskapsbudgeten och antalet gynnade områden .
jag tvingas i likhet med kollega mccarthy konstatera att antalet områden har skurits ned på ett ganska drastiskt sätt .
det vore önskvärt med en viss frihet för medlemsstaterna att inom en viss budget själva bestämma antalet projekt .
vad budgeten beträffar så består urban som sagt av stöd och komplettering till den nationella politiken .
om så behövs för att generera extra medel är det enligt min uppfattning också helt logiskt att i första hand vända sig till medlemsstaterna och privata finansiärer .
de gröna kan därför inte räkna med vårt stöd för ändringsförslag 2 , vilket de inte heller fick under utskottssammanträdet .
dessutom anser jag att stöd till en stad eller en trakt , i synnerhet där det handlar om gemenskapsbidrag , måste ha en stimulerande effekt .
strukturellt stöd skulle leda till bidragsberoende .
på det sättet skjuter vi över målet .
slutligen bara en allmän kommentar om interreg .
stöd till gränsöverskridande projekt skall enligt min uppfattning endast beviljas om regionerna verkligen önskar att få detta .
vid genomförandet av projekten är det också viktigt att de inte står i strid med den allmänna gemenskapslagstiftningen .
enligt revisionsrättens rapport för år 1998 är det inte någon inbillad risk .
det är också anledningen till vårt ändringsförslag för att förebygga motstridigheter mellan allmän politik och konkreta projekt .
jag tar mig friheten att först av allt uttrycka min bestörtning över de 14 rådsrepresentanternas förhastade fördömande av österrike .
herr talman , kära kolleger ! reformen av strukturfonderna leder till att gemenskapsinitiativen koncentreras till sammanlagt fyra .
jag välkomnar fortsättningen på och den framskjutna placeringen av interreg .
dock orsakar förseningen av direktivförslaget ett par problem .
regionerna inkluderades inte i tillräcklig utsträckning i förberedelserna till direktivet , trots att det under diskussionen om reformen av strukturformerna ofta krävdes att så skulle ske .
det saknas en direkt övergång mellan interreg ii och iii , vilket i praktiken drar med sig osäkerhet i planeringen och luckor i finansieringen .
det är synd , för det äventyrar verkligt meningsfulla projekt .
vid genomförandet av interreg måste samordningen och synkroniseringen med övriga berörda finansinstrument tryggas .
detta är särskilt viktigt för att höja effektiviteten av de beviljade anslagen .
problem uppstår dock särskilt i och med att anslagen beviljas årsvis och är knutna till projekt , exempelvis phare , i jämförelse med den flerårsbasis som gäller för interreg-anslag och det åtgärdsrelaterade anslagsbeviljandet .
detta kommer framdeles att medföra praktiska problem , men jag hoppas att det ändå blir möjligt att genomföra interreg på ett meningsfullt sätt .
herr talman , mina damer och herrar ! gemenskapsinitiativet leader har visat sig vara ett verktyg för att ge impulser till innovativ utveckling och till pilotprojekt i liksom från landsbygdsområdet .
därför är upprätthållandet av just detta gemenskapsinitiativ och den nya upplagan i leader + -programmet mycket välkomna .
det nya leader + -programmet kan nu tillämpas på hela landsbygdsområdet i europeiska unionen , vilket leder till bättre möjligheter för de projekt som skall stödjas .
det är viktigt att samordna leader + med övriga stödmöjligheter i europeiska unionen , men precis lika viktigt är det att samordna det med de andra nationella stöden .
det måste undvikas att stöden överlappar varandra , och samtidigt måste synergieffekter kunna utnyttjas .
i enlighet med detta måste målet att stärka integreringen av de olika leader-stödområdena verkligen välkomnas .
jordbruket är en av de bärande pelarna på landsbygdsområdet och måste kunna få del i leader-initiativet , eller också kan den strukturella förändringen i jordbruket få sällskap av leader-initiativet genom att nya arbetstillfällen skapas på landsbygden .
alla ekonomiska sammanhang som rör landsbruket måste uppmärksammas i leader + -programmet , och endast genom gemensamma ansträngningar kan man då nå det optimala .
leader måste nu förverkligas .
de operativa programmen måste beviljas av kommissionen så snart som möjligt , dvs. en praktiskt genomförd och effektiv hantering av förslagsställandet samt snabbast möjliga godkännande av förslaget .
fem månader har man räknat med .
det tycker jag är litet för lång tid .
man bör i detta fall försöka klara sig med kortare tidsfrister .
för den som har utvecklat ett projekt och fått det färdigt vill också sätta igång med genomförandet så snart det bara går .
trots all glädje över den nya utformningen av gemenskapsinitiativet leader + är det dock en sak som ligger mig varmt om hjärtat : europeiska kommissionen har i sitt förslag krävt ett övervakningscentrum för leader + -programmet utan att närmare gå in på hur förslaget skall genomföras .
detta innebär följande frågor för mig : vem skall arbeta där ?
hur väljs dessa personer ut ?
framför allt , varifrån kommer det kapital som behövs , och var skall detta övervakningscentrum vara beläget ?
jag menar nu att leader + -programmet inte behöver ett öre till ytterligare förvaltningsuppdrag , vilka det av naturliga skäl i alla fall skulle åligga kommissionen att utföra .
dessutom visar erfarenheten från andra områden där övervakningscentrer har inrättats att dessa förutom ett tvivelaktig skapande av nya arbetsplatser inte gör någon större nytta .
jag uppmanar därför kommissionen att själva och direkt sköta sina kontrolluppdrag samt att arbeta för en god utveckling av leader + -programmen .
dit hör ju också utvärderingen och offentliggörandet , vilket hittills ju också har varit fallet .
den största delen av de gränser som under sekler delat europa är tillskapade på ett konstlat sätt . de separerade unika geografiska områden och skapade starka skillnader i form av balanserad utveckling och sammanhållning .
våra inre gränser , eller det som är kvar av dem , ger inte längre upphov till krig , men de fortsätter att ge upphov till ekonomiska skillnader , sociala gränser och kulturell avskärmning mellan europas folk .
från gemenskapens institutioner måste vi arbeta för att komma över denna ärrbildning i gränsområdena , som är en motsättning till andan av europeisk enhet .
den ekonomiska och sociala sammanhållning som vi kämpar för konkretiseras genom interreg-initiativet , i den territoriella sammanhållningen och i integrationen av gränsområden och vår kontinents randområden .
interreg är sedan sin tillblivelse fröet till en verklig gemenskapspolitik för den fysiska planeringen av territoriet och en verklig polycentrisk uppfattning om det europeiska territoriet .
europaparlamentet beklagar bara att vi måste anta en resolution om detta initiativ , som vi håller med om , när vi ännu inte känner till utvärderingen av interreg ii .
men vi är medvetna om att det inte är lämpligt att dröja längre med tillämpningen av denna tredje utgåva , eftersom vi då skulle kunna riskera flera projekts framgång och en kontinuitet i de projekt som redan är igång .
interregs framgångar är uppenbara och det uttrycker de lokala , regionala och nationella myndigheter som deltagit i medfinansierade projekt .
att lära tillsammans , förnya , dela projekt och goda erfarenheter , förstå och tolerera varandra är några av de lektioner som deltagarna i detta initiativ kan lära av detsamma .
det finns en hel del intressanta frågor kring detta , observation , koncentrationsprincipen ...
jag skulle vilja uppehålla mig kring de förvaltande organen .
det är nödvändigt att söka gemensamma , interregionala och transnationella förvaltningsorgan i vilka alla lokala och regionala myndigheter deltar aktivt , samt de ekonomiska och sociala parterna .
parallella projekt på ena och andra sidan gränsen bör inte upprepas .
vi måste skapa en gränsöverskridande kultur och för detta ändamål är det nödvändigt att finna nya vägar när det gäller administrativt samarbete och med fantasi övervinna existerande hinder , samt övervinna de svårigheter de olika graderna av kompetens i varje medlemsstat , i varje region och i varje kommun innebär .
det får inte vara så att ett projekt inte kan genomföras på grund av samtalssvårigheter .
under diskussionerna i utskottet har vi också konstaterat svårigheten att samordna interreg med andra finansiella instrument av årlig eller tvåårig karaktär , som meda , tacis eller phare .
genom förslaget till resolution i parlamentet har man verkligen försökt uppmärksamma dessa svårigheter genom att formulera förslag till kommissionen som gör det möjligt att lösa dem och genom att uppställa rimliga tidsfrister för att genomföra nödvändiga ändringar .
herr talman ! mitt skäl till att bidra till denna debatt har att göra med att urban-initiativet - särskilt i irland - har varit mycket framgångsrikt och jag vill verkligen att europeiska unionen ger ytterligare bidrag på detta område .
det är ett tråkigt faktum att det finns flera hundra , om inte tusentals , samhällen i europeiska unionen som lider av en mycket allvarlig fattigdom och eftersatthet .
t.o.m. i medlemsstater och städer som är oerhört välmående finns det många som bor i getton , under levnadsbetingelser där det inte finns tillräckligt med moderna bekvämligheter , där utbildningen är bristfällig , där den fysiska infrastrukturen är underutvecklad och där narkotika och andra fenomen är mycket vanliga .
det verkar som om europeiska unionen , för att visa att den har en roll när det gäller att hjälpa europeiska unionens medborgare , måste hjälpa medlemsstaterna för att visa att unionen fungerar för dessa medborgare och deras familjer .
programmet har varit oerhört framgångsrikt i irland , på samma sätt som jag naturligtvis känner till att det varit framgångsrikt i andra länder .
det var litet långsamt under inledningsfasen här , men detta berodde på att det var nödvändigt att lokalbefolkningen själv utvecklade dessa program .
det är viktigt att de använder sin initiativkraft och sin egen kännedom om lokala förhållanden vid utvecklingen av detta initiativ .
det skulle vara mycket lätt att se till att få dessa program snabbt utvecklade och i rätt tid om man tog hjälp av externa sakkunniga , men detta skulle undergräva hela syftet med urban-programmet .
jag vill ta upp ytterligare en sak innan jag slutar : vi bör ställa krav på det sätt på vilket dessa medel tilldelas och den plats detta program utvecklas , i det avseendet att det sker i samband med en seriös urban-utvecklingspolitik .
detta är tyvärr inte fallet i irland .
jag applåderar det innovativa förhållningssättet inom equal-programmet och målet att få ut diskriminerade grupper på arbetsmarknaden .
utvecklingspartnerskapen är en mycket klok idé , trots att de befinner sig på experimentstadiet .
det finns emellertid framför allt två skäl till varför jag har betänkligheter rörande utvecklingspartnerskapen .
de borde vara tillgängliga för mindre grupper , tillgängliga i det avseendet att de skall kunna planera , genomföra och övervaka programmen .
vi måste ha ett stort mått av flexibilitet inom programmet .
jag har också innan uttryckt oro rörande användningen av jargong i stället för ett enkelt och tydligt språk , så att det blir tillgängligt för alla .
jag är glad att denna tanke godtogs i betänkandet , men jag kan inte stödja ändringsförslag 9 , eftersom detta ändringsförslag faktiskt inte alls skrivits på ett enkelt språk .
för det andra oroar det mig att vissa diskriminerade grupper har särskilda problem - t.ex. de handikappades situation i fråga om tillträde till sina arbetsplatser .
genom projekten bör man också särskilt ta itu med detta problem .
man bör titta på dessa frågor samtidigt som man fastställer programmen .
jag har sannerligen för avsikt att göra detta tillsammans med organisationer och grupper i min valkrets i west midlands .
låt mig nu ta upp den kontroversiella frågan om asylsökande och flyktingar .
även om jag inte stöder att de flyktingar som förvägrats flyktingstatus och hotats med avvisning skall få tillgång till equal-initiativet , stöder jag möjligheten till tillgång för alla övriga asylsökande och flyktingar .
det är bara rätt och riktigt att de skall kunna få tillgång till equal-initiativet på samma sätt som alla andra .
i betänkandet om leader är det landsbygdens utveckling som står i centrum .
det är inte så vanligt och det är därför glädjande , särskilt som leader-programmen varit huvudbeståndsdelar i unionens politik för landsbygdsutveckling .
det bör erinras om att dessa program inte bara varit strukturerande beståndsdelar för en politik för fysisk planering utan också grundläggande instrument för ekonomisk och social sammanhållning i områden som ofta är ömtåliga , exempelvis områden med utbredning av ödemark .
det är viktigt att betona att för att kunna komma i fråga för stöd enligt leader-programmet har de lokala aktörerna samarbetat , diskuterat och utarbetat projekt .
därför har dessa program varit viktiga för en demokrati där människor är delaktiga och för medborgartanken i europa .
konceptet leader + skall också innehålla alla positiva aspekter av tidigare program .
en viktig fråga uppstår alltså : varför skall vi efter att i tio år framgångsrikt ha bedrivit dessa program förpassa leader + till en experimentroll ?
finns det så många andra europeiska åtgärder som gör att man kan stoltsera med 800 originella specifika erfarenheter som varit ovanligt lyckade ?
hur länge tänker kommissionen fortsätta att behålla leader på experimentstadiet innan programmet tillåts ingå i det allmänna konceptet för landsbygdsutvecklingens mainstreaming ?
jag ställer mig också frågande till de minskade riktlinjer dit kommissionen vill förpassa leader + .
herr kommissionär ! när vi européer , efter seattle , kämpar för de många funktionerna i projekten för landsbygdsutveckling , varför då begränsas av kriterier med mycket otillräckliga medel ?
det är en miljöpartist som talar till er : försiktighetsprincipen och en hållbar utveckling kräver ett mycket mer varierat synsätt under många fler former .
i det sammanhanget föreslår kommissionen att vi ytterligare skall begränsa åtgärderna för samarbete med lokala aktionsgrupper till enbart kandidatländerna .
det skulle vara bättre , vilket också utskottet för regionalpolitik föreslår , att ha en förstärkt samordning mellan leader + och gemenskapens program för samarbete och partnerskap , såsom interreg , phare , sapard eller meda .
att vara solidarisk med östeuropa är nog bra , men det räcker inte .
traditionen från de tidigare programmen , med länderna i söder , särskilt kring medelhavet , får inte överges .
därför kan vi ännu en gång betona att det som saknas på jordbruksområdet och inom landsbygdsutvecklingen är medbeslutande , som skulle göra det möjligt för oss att verkligen få medel för att program som kräver samarbete och tvärgående åtgärder skulle kunna innebära framsteg .
herr talman ! jag har några mycket korta kommentarer .
vi diskuterar den nya programplaneringsperioden och de nya riktlinjerna för de fyra gemenskapsinitiativen , utan att ha tillgång till en egentlig och fullständig utvärdering av den föregående perioden .
det är mycket negativt .
programmen och målen är vanligtvis väldigt optimistiska , resultaten är emellertid inte alltid tillfredsställande , och ofta lämnar bristen på öppenhet i förening med projektens komplexitet stort utrymme för misshushållning och till och med bedrägerier .
de gemenskapsinitiativ som vi diskuterar kan under vissa omständigheter spela en positiv roll .
det är dock nödvändigt att de inte underställs mål och strävanden inom ramen för en mer allmänt negativ ekonomisk och social politik , utan att de utvecklar en egen , självständig roll .
till exempel innebär equal-initiativets anpassning till målen om anställbarhet och ökad elasticitet i förhållandet mellan arbetsmarknadens parter att det förvandlas till en ny version av de lokala sysselsättningspakterna .
utvidgningen av leader-initiativet till alla unionens områden innebär en risk för en ytterligare marginalisering av de mindre gynnade regionerna , till fördel för de mer utvecklade regionerna .
interreg-initiativet skall omfatta utvalda regioner , med särskilt betoning på randregioner , öregioner , bergs- och icke-bergsregioner , som till exempel artas län i grekland , som helt felaktigt har utelämnas i bilaga i till kommissionens meddelande .
herr talman ! detta parlament och kommissionen har bestämt att landsbygdsutveckling skall betraktas som ett prioriterat politikområde , och jag vill här i dag välkomna den ansvarige kommissionären , kommissionär fischler .
vår reaktion i samband med de stödbehov som finns på landsbygden har varit långsam , men jag antar att det är bättre sent än aldrig .
familjejordbruket har nu erkänts som ett viktigt inslag i den europeiska jordbruksmodellen och är ett mål som skall diskuteras inom ramen för agenda 2000 .
jag anser att det inom de kommande fem åren kommer att fattas beslut som bestämmer framtiden för tusentals familjejordbruk som befinner sig på marginalen .
det anstår oss alla att göra allt som står i vår makt för att säkerställa deras fortlevnad .
som kommissionären känner till kommer inte bara jordbruksnäringen att vara tillräcklig för att säkerställa en hållbar utveckling på landsbygden .
av detta skäl behöver vi en samordning av alla politikområden som kan spela en positiv roll för landsbygdens utveckling .
i detta avseende har leader etablerats som ett effektivt utvecklingsinitiativ .
det ger möjligheter för lokala samhällen att fastställa sin utvecklingspotential och att aktivt delta i en diskussion av dessa problem .
det frivilliga deltagandet i utvecklingsprogram är inte alltid något som uppskattas fullt ut .
genom leader kan det emellertid inte råda några tvivel rörande effektiviteten i detta sammanhang som en integrerad del av en bredare eu- och nationell politik .
samtidigt som jag sammanfattningsvis välkomnar godkännandet av leader + , oroas jag av tidsglappet mellan avslutandet av leader ii och inledningen av det nya programmet .
jag uppmanar er att ta allvarligt på detta problem .
ett avbrott i verksamheten kommer att få allvarliga konsekvenser för programmet och en störande effekt på de frivilliga och yrkesmässiga arbetsinsatserna .
herr talman , herr kommissionär , mina damer och herrar ! efter att ha fått kännedom om meddelandet från kommissionen om initiativet interreg iii , och med tanke på att jag inom ramen för utskottet för regionalpolitik , transport och turism deltagit i omröstningen om decourrières betänkande , vill jag inte bara uttryckligen säga att vi principiellt är överens dels om initiativet , såsom det föreligger , och särskilt inom ramen för interreg iii b , och dels om att kommissionen skall godkänna den verksamhet som bidrar till att återupprätta landskap som lidit skada på grund av jordbrukspriserna , en sektor där ett stort antal föreningar , särskilt på jaktområdet , redan gör enorma satsningar i mitt land .
jag vill också ge mitt uttryckliga stöd till kommentarerna från utskottet för regionalpolitik , transport och turism , framför allt när det gäller att beklaga bristen på integration av de yttersta randområdena inom område a i programmet , eller påpeka bristen på precision när det gäller urvalskriterierna för villkoren för genomförande av område iii c , och slutligen när det gäller att kräva att parlamentsledamöterna skall vara delaktiga i ett europeiskt övervakningscentrum för gränsöverskridande , transnationellt och interregionalt samarbete .
jag vill också uttrycka ett verkligt förbehåll mot tendensen i kommissionens meddelande att , enligt interreg iii och iii b , knyta miljöskyddet enbart till utvecklingen av natura 2000 , som förefaller mig ofta vara ett alltför abstrakt medel för att försvara de ekologiska system , vars användare riskerar att uteslutas eller starkt begränsas .
jag skulle avslutningsvis vilja betona , genom att i förväg be om förståelse från kommissionen och berörda ministerråd , att det skulle vara lämpligt att ytterligare informera de europeiska folkvalda om de förfaranden som är knutna till inrättandet av interreg-ärendena och liknande initiativ .
och vi måste dessutom ytterligare införliva dem i processen med att utarbeta och genomföra berörda program , annars blir det svårt att förstå och försvara deras roll mot lokala och nationella myndigheter och till och med mot medborgarna .
herr talman ! först och främst skulle jag vilja framföra ett hjärtligt tack till föredraganden för equal-betänkandet , stenzel , för allt som hon har gjort för att för att vi allesammans skall få insikt i detta svåra ärende .
equal är ett mycket svårt program eftersom man där försöker att sammanföra så många gamla program och ändå vill se över dem på ett nytt sätt , och detta med mindre pengar än vad som stod till förfogande i de tidigare fonderna .
det är bara antalet personer som berörs av dessa program som egentligen inte har minskat .
därför är det mycket svårt att få en balans till stånd , inte bara mellan de olika länderna , inte bara mellan de olika delarna , utan i synnerhet även mellan de olika grupper som nämns i programmet , och det är egentligen det som har sysselsatt oss fram till i dag .
här och där fälls kommentarer om att den ena gruppen måste få mer än den andra .
själv har jag särskilt ägnat mig åt de handikappades och de äldres ställning inom ramen för programmet , och jag måste säga att de handikappade och de äldre hade kunnat bli helt bortglömda om inte europaparlamentet hade ägnat sig åt den frågan så intensivt .
en del andra grupper har nämnts , men det är framför allt medlemsstaterna som ligger på lur .
jag känner till exempel till en medlemsstat som vill använda en stor del av hela programmet till en enda del , nämligen flyktingarna .
jag skulle därför vilja be kommissionären att ordentligt se till att det upprättas en balans mellan de olika grupperna .
det får inte vara så att en medlemsstat , genom att åberopa subsidiaritetsprincipen som förevändning , kan säga att allt skall gå till en enda grupp .
jag tror att det krävs sträng tillsyn i detta fall , för annars får man just det som meijer varnade så starkt för , nämligen att det kommer att uppstå etablerade intressen och att människor tänker att pengarna är deras .
det är inte på det sättet !
de måste varje gång fördelas på nytt .
det skall handla om innovativa projekt , och det får inte vara så att de helt och hållet försvinner in i finansministerns kassa .
det är inte syftet , och det är en viktig punkt som vi måste beakta här .
jag tror att de kvarvarande problem som vi har haft inom parlamentet , som till en stor del härstammar från det faktum att det är så svårt att göra denna avvägning , kan lösas .
vad kommissionen beträffar hoppas jag att den kommer att kunna ansluta sig till den kompromiss som kommer att nås här i parlamentet och som framför allt är inriktad på balans .
för att ytterligare understryka detta - situationen är naturligtvis aningen svår - har parlamentet för enkelhetens skull och för säkerhets skull tills vidare placerat equal-programmet i reserven , så att parlamentet så småningom skall bli övertygat om på vilket sätt genomförandet kan komma till stånd .
jag tror att det också är positivt .
parlamentets ställning i hela denna procedur är litet otydlig .
även i arbetsordningen är denna ställning otydlig , och just därför är det mycket bra med denna reserv .
värderade kolleger ! det är ett oemotsägligt faktum att interreg-initiativet stöder ansträngningarna att nå ekonomisk och social sammanhållning i europeiska unionen .
jag vill dock betona den särskilda betydelse som interreg har för balkanregionen , där de senaste årens politiska utveckling och krigshandlingar har fått stora ekonomiska konsekvenser för grannländerna , särskilt för mitt land , grekland , som är det enda medlemslandet som är beläget på den hårt drabbade halvön .
för grekland , grannländerna italien och österrike , men även för hela europa , är balkans sociala och ekonomiska återuppbyggnad , som skall leda till politisk stabilitet , en fråga av största betydelse .
fram till i dag har vissa av länderna på balkan fått stöd genom phare- och obnova-programmen , andra inte .
under den nya programplaneringsperioden , inför utvidgningen och med hänsyn tagen till att stöd genom nya stödinstrument och förordningar , som till exempel ispa och sapard har planerats , är det absolut nödvändigt att samordna stödet på interregs tre insatsområden med det övriga stödet till tredje land .
vi välkomnar följaktligen formuleringarna om detta i kapitel 7 i europeiska unionens text om fastställande av interreg-riktlinjer .
ansträngningarna för att samordna och följaktligen effektivisera planeringen måste fördelas lika på alla program , och jag säger detta eftersom det i meda-programmet , under den föregående perioden , fanns vissa problem som bör lösas , så att vi behandlar alla de tredje länder som deltar i programmet lika .
jag skulle vilja avsluta , herr talman , med att konstatera att man i den nya planeringen av områdena för mellanstatligt samarbete inte har tagit hänsyn till medelhavsområdets geografiska egenhet , som borde rättfärdiga skapandet av ett särskilt område för kust- och öregioner .
vi begär alltså av kommissionen att den särskilt skall beakta frågan om samarbete i havsnära regioner och i öregioner vid kommande revideringar av områdesplaneringen .
avslutningsvis , herr talman , betonar jag nödvändigheten av att europeiska unionen insisterar på denna slags initiativ , som avser att utplåna orättvisor mellan våra regioner och att få till stånd en harmonisk utveckling för dem .
och eftersom det i dag är alla hjärtans dag , föreslår jag , som gammal borgmästare i en regional stad , att vi alla förklarar vår kärlek till de europeiska regionerna , de som behöver den kärleken .
herr talman ! jag vill tala om equal-betänkandet , särskilt frågan om flyktingpolitik .
i förra veckan diskuterade vi den österrikiska regeringsbildningen med stort engagemang .
i dag diskuterar vi redan den österrikiska regeringskoalitionens flyktingpolitik , eftersom stenzel som har författat equal-betänkandet ju representerar det österrikiska konservativa regeringspartiet och dess politik .
det mest uppseendeväckande i hennes ursprungliga betänkande var att hon ville begränsa flyktingstödet till den lilla grupp flyktingar som omfattas av genèvekonventionen , dvs. så kallade kvotflyktingar eller fn-flyktingar .
i själva verket är det de andra flyktingarna , nämligen de som står utanför kvoten och fn-stöd , som har det största behovet av stöd .
utskottet förkastade detta diskrimineringsförslag och beslutade att alla flyktingar skall få plats i equal-programmet på lika villkor .
en del av utskottet solidariserade sig emellertid med stenzels förslag och formuleringar .
det betyder enligt mitt sätt att se att haiderpolitiken redan kastar sin skugga över detta parlament .
därför är det av avgörande betydelse att kammaren med största möjliga eftertryck slår fast att alla flyktingar skall ha plats i equal-programmet .
jag vill till sist säga att jag hade vissa betänkligheter i förra veckan när vi diskuterade regeringsbildningen , men när det gäller att diskutera och kritisera den österrikiska flyktingpolitiken , då har jag inga betänkligheter .
jag hoppas att engagemanget i kammaren blir lika stort denna gång .
herr talman ! under eu : s senaste budgetplan från 1994 till 1999 , när det fanns 13 olika initiativ i kraft , var det gränsöverskridande interreg ii-programmet ett viktigt initiativ .
det faktum att nästa strukturfondsrunda mellan 2000 och 2006 omfattar interreg-initiativet anser jag vara en mycket tydlig fingervisning om den betydelse som tillmäts detta av eu : s medlemsstater .
interreg i-programmet mellan 1989 och 1993 och interreg ii-programmet mellan 1994 och 1999 har visat sig vara en fullständig framgång när det gällt att skapa ett närmare samarbete mellan angränsande medlemsstater i frågor som rör social och ekonomisk utveckling .
eftersom jag själv kommer från gränstrakterna i nordvästra irland har jag sett den viktiga roll som interreg i och ii har spelat under årens lopp , och jag är glad att kunna välkomna interreg iii .
kommissionen kommer att tilldela 67 miljoner pund till interreg iii-programmet , som kommer att användas till en fortsatt utveckling av gränsöverskridande ekonomiska projekt mellan irland och nordirland .
europeiska unionen har spelat en viktig roll vid utvecklandet av gränsregionerna i irland under årens lopp .
europeiska unionen är den enskilt största bidragsgivaren med 80 miljoner pund till internationella fonden för irland .
europeiska unionen bidrar med 75 procent av det totala freds- och försoningsprogrammet .
sammanfattningsvis har interreg , internationella fonden för irland och freds- och försoningsprogrammet spelat en viktig roll för den löpande fredsprocessen .
herr talman ! jag skall tala om interreg och bland annat för att respektera tidsbegränsningen hålla mig till några få kritiska punkter .
vi har alla gett uttryck för en positiv syn på att detta program förlängs och på utvidgningen av insatsområdena till att förutom samarbete över gränserna även omfatta samarbete mellan nationer och regioner .
detta hindrar dock inte att vi är medvetna om det faktum att större delen av resurserna - mellan 50 och 80 procent - kommer att reserveras för samarbetet över gränserna , för volet a i interreg iii-programmet .
det val man sedan har gjort , att för detta volet befästa de nuvarande samarbetsområdena , vad gäller vilka regioner som äger tillträde , anser vi fortfarande är både felaktigt och motsägelsefullt .
vi hoppas verkligen att kommissionen kommer att se över detta och vidgå parlamentets ståndpunkt i sak , och inte som en formell aktningsbetygelse .
samarbetet över gränserna sker fortfarande nästan uteslutande över landgränserna och på de ställen man har gjort undantag för vattengränser saknas insyn i besluten och de bär ofta spår av kompensation för andra delar av gemenskapspolitiken .
diskrimineringen framstår som enormt mycket allvarligare för öarna , vilkas regionala förhållanden inte kan annat än präglas av att de uteslutande har havsgränser .
detta är i linje med en diskriminering som man fortsätter att tillämpa utan att ta hänsyn till artikel 158 i fördraget , som gäller öregionerna i sammanhållningspolitiken .
det är ännu mer allvarligt att detta sker utan hänsyn till den nya väg vi har slagit in på i och med utvidgningen till regioner som malta .
härav de förslag vi har lagt att utvidga de regioner som kan komma i fråga åtminstone till siciliens nuts iii-gränser gentemot malta och för alla de adriatiska regionerna gentemot balkan .
herr talman , herr kommissionär , kära kolleger ! jag skulle vilja uttrycka min tacksamhet över att kunna konstatera att de yttersta randområdena , däribland de franska utomeuropeiska departementen , varit föremål för ett visst intresse inom ramen för initiativet interreg iii , vilket öppnar nya perspektiv för att de skall kunna samarbeta med länderna inom sitt geografiska område , även om man kunde ha hoppats på något bättre , bl a när det gäller tillgång till de olika områdena .
under lång tid har våra regioner haft blicken fästad på sin europeiska huvudstad , sannolikt en kvarleva från kolonialtiden , och struntat i och till och med föraktat sina närmaste grannar .
detta hör i dag absolut till det förgångna .
våra regioner har blivit medvetna om att de tillhör en miljö som de är knutna till , inte bara geografiskt utan också genom sin kultur och sitt folks historia , vilket ger upphov till en stark strävan efter en djupare förankring i denna miljö .
men denna insikt handlar inte bara om identitet .
den är också beroende av en rättvis uppskattning av våra tillgångar .
la réunion befinner sig exempelvis mitt i axeln för utbyte mellan länderna i södra afrika och de i sydostasien .
ön kan inte stå vid sidan om de regionala grupperingar som verkar i området , eftersom den då riskerar att gå miste om en historisk möjlighet , och detsamma gäller våra regioner i västindien .
avslutningsvis är vi övertygade om att våra ungdomar kan skönja en utväg ur den dramatiska arbetslösheten som gör dem förtvivlade , om vi till intilliggande länder kan exportera den know-how som förvärvas tack vare strukturfondernas åtgärder .
utnyttjandet av interregs anslag kan göra våra regioner till verkliga brohuvuden för europeiska unionen inom deras geografiska områden , och på så sätt ge dem en världsomspännande dimension .
jag räknar med kommissionen och särskilt med er , herr kommissionär , för att ge dem medel till effektiva åtgärder .
herr talman , kommissionärer ! jag välkomnar varmt möjligheterna till ett ökat europeiskt samarbete i samband med interreg , men jag oroar mig för att förslaget ger färre möjligheter för havsområdena än för andra områden i detta avseende .
jag förstår kommissionens egen oro över att geografiskt avstånd kan inverka menligt på ett effektivt samarbete .
det finns i vilket fall många havsområden som redan upprättat kontakter .
olika lokala myndigheter i nordsjöområdet är ett bra exempel på detta .
interreg skulle mycket väl kunna förstärka detta samarbete .
som ett resultat av detta vill jag se att det görs vissa mindre ändringar av riktlinjerna för att skapa litet mer flexibilitet och för att anpassa de sätt på vilka havsområdenas intressen kan hamna mellan område a och område b. dessa anpassningar omfattar ett förtydligande av möjligheterna för samarbete mellan havsområden och tillåtande av en bredare utveckling av praktiska och genomförbara projekt , i synnerhet de som har en infrastrukturell karaktär .
sådana åtgärder kommer att likställa havs- och öområden med andra områden i eu .
jag hoppas att de blir antagna .
herr talman ! vår grupp välkomnar den övergripande kraften hos equal-initiativet genom att , om du är en brittisk muslim som har någon form av fysiskt handikapp inte längre behöver välja mellan vilken diskrimineringskategori man tillhör som målgrupp : man kan använda sin sakkunskap och erfarenhet för att lösa problem , i stället för att betraktas som själva problemet .
det finns mycket sakkunskap inom de relevanta organisationerna som är värd att dela med sig av .
vi välkomnar också erkännandet av behovet av utvärdering och spridning av bästa metoder för åtstramning av den gränsöverskridande nivån .
vi är därför bekymrade över , som andra har nämnt , antalet ändringsförslag som försöker att ytterligare marginalisera en del av de i samhället som redan tillhör de mest marginaliserade , genom att förespråka en mycket snäv definition av &quot; flykting &quot; .
min grupp kommer inte att stödja dessa ändringsförslag .
vi är också bekymrade över det antal ändringsförslag som innebär att man genom att försöka införa en större flexibilitet , kanske löper en risk att skapa förvirring när det gäller var ansvaret för equal-initiativets verksamhet ligger .
herr talman ! det gläder mig att se att urban-initiativet ges en mer helhetlig inriktning och att man med initiativet försöker lösa sammanhängande problem .
det finns dock , herr talman , en risk med denna utspridning : att våra försök att uppfylla många mål leder till en övergripande ineffektivitet .
varje enskilt fall av tillbakagång i ett stadsområde är naturligtvis speciellt .
det finns emellertid en resultant , en hård kärna , som består i att arbetslösheten ökar , att de offentliga tjänsterna försvinner eller skärs ned samt att små och medelstora företag , affärer och andra inrättningar försvinner .
jag skulle önska att man med urban-initiativet först och främst riktade in sig på att försöka finna svar på dessa orsaker till tillbakagång i städerna .
och då är det naturligtvis nödvändigt att nå samförstånd och att samordna den centrala politiken med utvecklingspolitiken , så att även denna ges en ny inriktning och samverkar med målen i de urban-initiativ som genomförs i våra länder , i stället för att helt enkelt lägga fram de där programmen som ett alibi för frånvaron av en sådan politik .
herr talman , herr kommissionär , kära kolleger ! jag begränsar mitt inlägg till francis decourrières betänkande .
programmet för gemenskapsinitiativet interreg är ett extremt viktigt verktyg när det gäller europeisk utveckling och fysisk planering , särskilt om vi effektivt skall beakta förhållandet mellan europeiska unionens centrum och dess randområden .
interreg skall därför vara ett instrument som främjar unionens territoriella sammanhållning , om vi vill undvika ett europeiskt territorium uppdelat i två eller tre hastigheter .
det förefaller mig självklart att de regionala och lokala myndigheterna , de organisationer som företräder dem , regionkommittén och självfallet europaparlamentet , tydligare och så snart som möjligt skulle ha kopplats in när det gäller att utarbeta programmet .
men man måste konstatera att så inte var fallet när kommissionen förberedde sitt meddelande , som offentliggjordes den 13 oktober förra året .
även om jag godkänner de allmänna riktlinjerna för interreg iii , förefaller det mig ytterligt viktigt att se till att det finns en bättre förbindelse mellan detta program - som finansieras av europeiska regionala utvecklingsfonden ( eruf ) - och övriga fonder för yttre samarbete , däribland bl.a. europeiska utvecklingsfonden avsedd för avs-länderna .
i det hänseendet skulle jag vilja tacka utskottet för regionalpolitik , transport och turism för att ha antagit ett av mina ändringsförslag som lägger till europeiska utvecklingsfonden ( euf ) i förteckningen över dessa fonder .
de yttersta randområdena , bl a de fyra franska utomeuropeiska departementen , måste kunna samordna interreg iii och euf för att också de skall kunna finansiera samarbetsprojekt med sina avs-grannar inom respektive geografiska område .
jag ber också kommissionen att vänligen på nytt överväga de dåliga möjligheter som erbjudits de yttersta randområdena och öregionerna enligt riktlinjerna i meddelandet .
dessa regioner skall , liksom samtliga övriga regioner i unionen , kunna utnyttja interreg iii fullt ut , särskilt som programmet regis , som var avsett för dem , nu avskaffats .
avslutningsvis vill jag beklaga de låga ekonomiska bidrag som avsatts för område c , avsett för samarbete mellan regioner , och vars betydelse inom gemenskapen ändå inte kan förnekas .
herr talman ! min utgångspunkt är equal-betänkandet och jämställdhet mellan män och kvinnor , även om jag måste erkänna att det emellanåt är tröttsamt att tala om denna fråga som har fått upprepandets natur , i varje fall när man är i min ålder .
men det är tyvärr nödvändigt att återigen påpeka att vi inte uppnått jämställdhet .
men kanske kan ett genombrott här leda fram till ändringar på andra områden .
för mig betyder nämligen inte jämställdhet att båda parter i ett äktenskap arbetar hela tiden och lämnar barnen till en dagmamma , dvs. en invandrare , som inte har fått en chans att få ett annat jobb .
om det skall vara så har vi inte kommit någonvart sedan solkungarnas tid .
nej , jämställdhet innebär att vi alla deltar i både arbetslivet och familjelivet .
utvecklingen går tyvärr inte i den riktningen , tvärtom .
jag tycker därför att punkt 7 innehåller något mycket viktigt .
här står nämligen : &quot; equal kommer att användas som försökslaboratorium för utveckling och förmedling av nya metoder för genomförande av sysselsättningspolitik &quot; .
man får hoppas att det lyckas .
herr talman ! i samband med arbetsordningen vill jag bara säga att om jag inte är här när kommissionen svarar - inte därför att jag ställt några särskilda frågor , men jag hoppas dock att kommissionen har gjort efterforskningar - beror detta på att det samtidigt med denna debatt pågår ett sammanträde i utskottet för kvinnors rättigheter och jämställdhetsfrågor om kvinnor i beslutsprocessen .
herr talman , mina damer och herrar ! de som ägnar sig åt landsbygdsområdet vet att leader-programmet , såväl leader i som leader ii - och jag hoppas även leader + - hör till berättelserna om de framgångar som europeiska unionen har lanserat .
framgångarna kom sig även av att leader-programmens grundkoncept framkallade en mycket stor aktivitet hos den berörda befolkningen .
det gläder mig att grundsatsen för leader + har stannat vid detta grundkoncept .
det finns dock ett problem som vi måste ta itu med gemensamt .
eftersom leader är något som kan liknas vid en verkstad med ett bottom-up-koncept , är det enormt många idéer som under årens lopp har mognat genom leader i och ii , idéer som så småningom förstås inte är så helt nya och framgångsrika längre .
och på grund av framgångarna leder grundsatsen naturligtvis till att de en vacker dag faller bort ur leader .
därför måste vi se till att det som har visat sig vara framstående i de bra leader-projekten inte plötsligt avbryts , utan de idéer som har visat sig vara goda någon gång måste föras över till de normala programmen som en fast , positiv komponent i stödet till landsbygdsområdet .
det är ju också grundidén .
att genom nya idéer i leader prova något , tillsammans med de inblandade på plats , med de kommunala sammanslutningarna på plats , med många oberoende organisationer , med kyrkorna , tillsammans med alla som har hjälpt till att verkligen få igång nya idéer på landsbygden .
här måste vi se till att de positiva saker som verkligen sticker ut på något sätt blir en fast beståndsdel i ett förnuftigt arbete inom landsbygdspolitiken .
nu ber jag kommissionen : ge akt på att de organisationer och de befolkningsdelar som satsar sin kompetens också verkligen tas emot .
det får inte vara så att man försöker sig på att mer eller mindre marginalisera den eller den organisationen som bildas just för att bidra med en ny idé och som ännu inte är särskilt känd - och må det så vara på grund av officiell politik på lokal eller regional nivå .
stanna kvar vid de positiva erfarenheter som leader hittills har visat .
i början kan det ibland vara litet som att lägga ut rökridåer att säga att det är för idealistiskt uttänkt .
och sedan under arbetets gång , under genomförandet , framträder det så småningom något som den officiella politiken - även vi på vår nivå - inte alls kunde föreställa sig , att det plötsligt skulle mogna och bli så bra .
det är detta som har varit charmen med leader , och det får bara inte gå förlorat !
herr talman ! jag välkomnar equal-initiativet och betänkandet i vilket man betonar behovet av att skilja mellan åtgärder för bekämpning av diskriminering av kvinnor och åtgärder för bekämpning av diskriminering av minoritetsgrupper .
kvinnor tillhör ingen minoritet och kvinnor drabbas ofta av dubbel diskriminering som medlemmar av minoritetsgrupper , såväl som på grund av sitt kön .
detta är skälet till varför det behövs särskilda åtgärder för kvinnor , såväl som mainstreaming .
detta tas upp i betänkandet och man föreslår en integrering av åtgärder för att åstadkomma jämlikhet mellan kvinnor och män i alla arbetsaspekter ; man tar också upp betydelsen av samarbete med de lokala och regionala organ som finns närmast medborgarna , för att se till att alla projektresultat har granskats ur ett jämlikhetsperspektiv .
deltagandet av frivillig- och gemenskapsgrupper kommer också att bli en viktig del av equal-initiativet och projekten .
utvecklingspartnerskapen inom ämnesområdena , vilka anges i ändringsförslag 22 , skulle göra det möjligt även för de mindre organisationerna att spela en roll inom equal-initiativet .
min grupp kommer att stödja ändringsförslag 22 .
herr talman , ledamöter ! det betänkande kammaren diskuterar i dag är otvivelaktigt mycket viktigt .
styrkan i gemenskapsinitiativet interreg för programplaneringsperioden 2000-2006 är , förutom de mål det syftar till , det mervärde det innebär i ljuset av den numera snart förestående utvidgningen av europeiska unionen till att omfatta nya länder i östeuropa och medelhavsområdet .
det är just inför denna händelse som europeiska unionen enligt min mening måste ta krafttag för att minska de regionala skillnaderna och sätta stopp för gränsområdenas isolering .
de sistnämnda har faktiskt - det bör man komma ihåg - en viktig roll att spela : rollen som broregioner gentemot de kandidatländer som kommer att bli medlemmar i unionen .
det är just mot bakgrund av detta som jag har lagt fram några ändringsförslag som jag anser är ytterst viktiga och som utskottet för regionalpolitik , transport och turism har gjort till sina .
med dessa vill vi utöka de områden som kan komma i fråga för samarbete över gränserna till alla adriatiska regioner liksom de sicilianska provinser som har gräns mot malta - kandidatland i utvidgningen - vilka i dag oförklarligt nog inte omfattas av avsnitt a i bilaga 1 .
jag förlitar mig på att kommissionär barnier och europeiska kommissionens ordförande tar vederbörlig hänsyn till parlamentets ståndpunkt i frågan , i enlighet med uppförandekoden .
det är ett grundläggande intresse för hela europa att främja samarbete med kandidatländerna och ingripa till stöd för gränsregionerna .
slutligen anser jag att det är önskvärt att man söker förbättra samordningen mellan interreg-initiativet och de redan befintliga gemenskapsprogrammen som har extern politisk bärighet för bättre integrering och samordnad behandling av programmen .
herr talman , herrar kommissionärer , kära kolleger ! leader i var en verklig framgång , framför allt tack vare den flexibla administrativa förvaltningen mellan kommissionen och de lokala aktörerna .
jag tycker att det är beklagligt att kommissionen inte upprättat samma bokslut över leader ii , ett bokslut över projektens kvalitet , mängden förbrukade anslag och framför allt över att vissa lokala aktörer givit upp inför den administrativa och ekonomiska tungroddhet man stött på .
jag gläds emellertid åt att nya medel inrättats , inom ramen för leader + , för att hjälpa landsbygdsområdena att utveckla sin potential och genomföra målsättningarna med lokal och hållbar utveckling .
jag vill särskilt betona experiment med nya former för att förädla natur- och kulturarvet och förstärka den ekonomiska miljön , för att främja sysselsättningen .
jag tror man kan anta att utbyte av dessa positiva erfarenheter av utvecklingen också kan förekomma inom ramen för det gränsöverskridande samarbetet .
det är också intressant att notera att alla landsbygdsområden är stödberättigade enligt leader ii .
om emellertid möjligheten kvarstår för medlemsstaterna att , inom ramen för detta initiativ , fastställa områden , bör kommissionen se till att det finns en viss koncentration av resurserna och prioritera projekt inom mindre framgångsrika områden .
det krävs naturligtvis öppenhet om urvalskriterierna när det gäller projekt och lokala aktionsgrupper .
det förefaller mig också som om man framför allt skulle behöva se till att staternas eller de lokala myndigheternas ekonomiska system inte längre är de som orsakar betalningsförseningar , något som försatt vissa lokala aktionsgrupper i konkurs inom ramen för leader ii .
herr talman ! som ledamot från ett yttre randområde måste jag säga att det är en mycket speciell eftermiddag när det gäller regionalpolitiken och det säger jag med anledning av debatten om två gemenskapsinitiativ , urban och interreg .
jag vill påminna om att nämnda initiativ syftar till att , när det gäller det första , urban , att förbättra livskvalitén för medborgare som bor i stadsdelar i olika europeiska städer , och interreg , att främja sammanhållningen och att se regionernas mångfald och möjligheter i europeiska unionen , särskilt när det gäller att inkludera de yttre randområdena i kapitel b och c.
vi beklagar , precis som föredraganden , att kapitel iiia har tagits bort .
vi anser att hänvisningen i interreg att skapa ett europeiskt övervakningscentrum om samarbetets effekter är mycket klokt .
tack till föredragandena , särskilt decourrière för hans känslighet för de regionala frågorna och för att han accepterat våra ändringsförslag .
jag hoppas att kommissionären godkänner det förslag vi lägger fram .
herr talman ! när det gäller de olika initiativ vi behandlar denna eftermiddag vill jag strikt uppehålla mig kring en reflektion kring ett av dessa .
det gäller rent konkret urban-programmet . det är sant att vi i dag debatterar detta program eftersom europaparlamentet envisades med att det skulle vara kvar .
kommissionens förslag var att ta bort det , tillsammans med andra initiativ , men parlamentets förslag och kommissionens egen känslighet när det kom till kritan gjorde att urban-programmet bibehålls .
jag tycker att vi skall glädja oss över det .
men , vilka var kommissionens argument , och i synnerhet kommissionär monika wulf-mathies samt generaldirektör eneko landaburu , för att urban-programmet inte skulle vara kvar ?
argumentet var tungt .
den urbana frågan är så viktig att vi inte kan begränsa den och nästan nedvärdera den med ett program som har en väldigt liten budget .
i dag har vi programmet och jag tror således att vi uppnått något viktigt , detta tecken på identitet som urban är för europeiska unionen .
men jag skulle vilja vända mig till kommissionär barnier för att lägga vikt vid kommissionärens och generaldirektörens argumentation eftersom jag tror att de hade väldigt rätt .
den urbana dimensionen bör innefattas oerhört mycket djupare i alla strukturfonder .
den budgetnivå våra städer behöver - där 80 procent av den europeiska befolkningen lever och som till stor del håller på att utvecklas till det goda och det dåliga vi har i europa - , tror jag kräver att denna europeiska dimension beaktas och urban-programmet får inte vara rättfärdigandet för att inte på djupet analysera , att inte prioritera och därför inte införa ett budgetanslag som vida överstiger det tidigare i program som påverkar städerna genom alla de europeiska fonderna .
därför anser jag att det är onödigt att åter upprepa det antal faktorer som kräver denna investering i de urbana områdena , faktorer som är på dagordningen . jag skulle vilja förmedla till kommissionären att vi hoppas på förståelse för detta .
samtidigt som vi välkomnar det sektorsövergripande förhållningssättet som finns i det nya equal-initiativet , är det mycket viktigt att programmet behandlar de typiska former av diskriminering som i synnerhet skadar handikappade personer : fysiska hinder på arbetsplatsen som påverkar dem med begränsad rörlighet , visuella informationssystem som inte är till nytta för blinda anställda , arbetssystem som effektivt hindrar dem som har inlärningsproblem eller psykiska problem .
handikapporganisationer och handikappade personers icke-handikappade företrädare måste få lämplig insyn vid beslutsfattandets alla stadier .
detta är skälet till varför detta parlament har lagt fram punkterna 10 och 15 i resolutionen för att se till att medlemsstaterna inte skall kunna bortse från någon målgrupp .
de handikappade har alltför ofta uteslutits från listan .
eftersom handikappade inte utgör en enda homogen grupp - många döva ser t.ex. sig själva som en språklig minoritet som inte erhåller respekt för sitt eget språk och sin egen kultur - är det nödvändigt , vilket uttrycks i punkt 9 , att tillåta att vissa partnerskap bestäms som är specifika för ett särskilt handikapp eller en annan grupp .
equal-initiativet är fortfarande mycket viktigt också i regioner som min hemregion i östra england , som i princip inte kan komma i fråga för stöd från mål 1-fonderna . vi har haft extra starka incitament för att erhålla medel från gemenskapsinitiativ och kan uppvisa en utmärkt historik .
före detta adapt-projekt som sträcker sig från core-projektet - genom vilket man har utvecklat nya leverantörskedjor inom bilindustrin i bedfordshire - till standardhöjande projekt för mindre företag i hertfordshire i essex .
vi har sett hur now-projektet har hjälpt 70 kvinnor att få arbete i suffolk , av vilka många kunde komma och dela med sig av sina erfarenheter direkt med oss i europaparlamentet i bryssel .
equal-initiativet är fortfarande viktigt för oss , eftersom det är just i relativt sett mer välmående regioner där icke-kvalificerade arbetstillfällen försvinner , och det är denna typ av arbeten som kan vara en viktig första hållplats för dem som är diskriminerade på arbetsmarknaden .
till sist några ord om interreg .
egentligen är det rent nonsens att partnerskap som upprättats 1994 nu förlängs med undantag av nya interregionala förbindelser .
under denna period har hamnarna great yarmouth och harwich på essex-suffolk-norfolkkusten infört betydelsefulla nya transport- och ekonomiska förbindelser med partner i nederländerna .
jag uppmanar parlamentet att stödja vårt ändringsförslag 2 , vilket kommer att säkerställa flexibilitet genom att inkludera nya områden , i synnerhet när det gäller havsgränser .
herr talman , ärade kommission , ärade damer och herrar ! herr talman , jag vill för allas information komma med ett klarläggande .
förbundskansler schüssels regering fortsätter driva förre förbundskansler klimas socialdemokratiska regerings flyktingpolitik .
det förekommer ingen ändring av flyktingpolitiken i österrike !
landsbygdsområdena utgör över 80 procent av eu : s yta , och 25 procent av befolkningen lever här .
som bondkvinna och ledamot har jag alltid varit angelägen om att inte se jordbruket som något för sig , utan att se till hela landsbygdsområdet .
särskilt värdesätter jag en integrerad satsning på landsbygdens utveckling eftersom jag är övertygad om att man kan skapa en aktiv och attraktiv livsyta för alla endast genom att sammanföra alla yrkesgrupper och alla människor på landsbygdsområdet till en gemenskap , kort och gott - landsbygdsområdets mångfaldiga funktion .
det nya leader + -programmet hälsar jag särskilt välkommet på grund av dess omfattande karaktär .
det kommer i framtiden att bli möjligt att ha program inte bara i de enskilda stödområdena , utan i alla regioner inom eu .
denna horisontella satsning är vettig i och med att programmen för landsbygdens utveckling också är utformade så .
finansieringen kommer framdeles inte längre att skötas via tre fonder , utan då endast ur europeiska utvecklings- och garantifonden för jordbruket ( eugfj ) .
därför kommer det att krävas en höjning av kvalitén på programmen , för eugfj skall vara ett verksamt finansieringsinstrument .
högre precision vid urvalet kommer att leda till höjd effektivitet , för pengarna skall inte slösas bort planlöst .
jag vill också peka särskilt på den punkt som bildar en ansats till en integrerad och miljöanpassad utvecklingsstrategi .
detta innebär att det finns en stor sysselsättningspotential för framtiden på landsbygdsområdet , och vi måste utnyttja detta om vi vill ge människorna på landsbygden ett perspektiv .
därför är politik på landsbygden mer än politik bara för bönderna .
leader + skall komplettera redan befintliga program , undvika överlappning och dubbelfinansiering och bidra till en så omfattande utveckling som möjligt .
på så sätt kan leader + tillsammans med programmen i förordning 1257 / 99 backa upp andra stöttepelaren i den gemensamma jordbrukspolitiken ännu mer och åstadkomma bästa möjliga resultat för det samlade landsbygdsområdet .
herr talman , bästa kolleger ! jag är inte alltid stolt över vad det här parlamentet sysslar med , men urban-programmet är ett av de bästa exemplen på vår verksamhet , det uppstod just på parlamentets initiativ .
kommissionen ville avskaffa urban , men den här gången drog parlamentet det längsta strået .
det är bra att urban fortsätter , ty man har på lokal nivå fått goda resultat av det .
problemen i europeiska stadsområden håller på att bli värre ; som tur är delar vi nu åsikt med kommissionen .
majoriteten av europas befolkning bor i städer , deras problem är bland de viktigaste inom regionalpolitiken och mycket komplicerade frågor .
risken för utslagning är stor .
i många franska och engelska städer finns redan slumområden där många onda ting föds .
ingen av oss vill ha sydamerikanska favelas i europa .
vi måste agera nu innan det är för sent .
städerna spelar också en avgörande roll för den europeiska ekonomin .
vi återkommer alltid till samma europeiska grundproblem : vårt näringsliv är inte tillräckligt dynamiskt och uppmuntrar inte individen i tillräckligt hög grad .
näringslivet måste vara starkt om vi skall kunna ta hand om våra närstående och vår miljö .
detta är inte politik utan livets enkla logik .
när det gäller användningen av pengar är det bra att pengarna nu har centraliserats , ty om man sprider skotten åt alla håll försvinner krutet all världens väg som en flock sparvar .
nu måste vi koncentrera oss på att lösa de små och medelstora städernas problem eftersom de inte har tillräckligt med kritisk massa .
på det sättet kan vi också ge mera fart åt de omgivande landsbygdsregionerna ; man glömmer ofta att städernas och landsbygdens problem i själva verket går hand i hand .
grunden för allt är att man skall uppmuntra individens innovativa förmåga och företagsamhet eftersom den massrörelse som skapar en intern regional reform börjar hos en individ .
att ge finansiering utan att det finns en ekonomi som står på egna ben är som att bära vatten till en sinad brunn : drickat räcker för en stund , men i morgon är brunnen åter tom.
herr talman ! i och med att interreg iii förverkligas går den europeiska samarbetspolitiken in i en ny fas .
vår uppmärksamhet riktas inte längre enbart mot de inre gränserna , utan även mot de yttre .
i dagens läge med globalisering och kulturell öppenhet behöver europeiska unionen instrument för att stärka sina band och sina kommunikationskanaler med angränsande regioner , särskilt i öst- och sydeuropa .
unionens gränser får inte längre utgöra ett hinder för en balanserad utveckling utan tvärtom en möjlighet , en bro till ett mer fruktbart samarbete .
via de ändringsförslag som har antagits i utskottet försöker parlamentet komplettera kommissionens arbete genom att föra in nya namn på listan över mottagarområden för stöden , särskilt till förmån för de yttre havsgränserna i sydeuropa .
i sitt förslag till riktlinjer påpekar kommissionen faktiskt att dessa gränser fordrar större uppmärksamhet än tidigare .
detta med beaktande av utvidgningsprocessen mot öst och processen för större integrering med medelhavsländerna .
som ordförande prodi också påminde om när han lade fram de strategiska målen för 2000-2005 är nylanseringen av barcelonaprocessen en prioriterad fråga för unionen , och interreg iii-initiativet kan ge sitt bidrag till att detta strategiska mål uppnås .
vi gläder oss åt det utmärkta arbete föredraganden har gjort och hoppas bara att kommissionen tar vederbörlig hänsyn till de förslag parlamentet har lagt fram , i enlighet med åtagandena i uppförandekoden för genomförande av strukturpolitik , och med de ändringar som behövs bekräftar detta gemenskapsinitiativs omvandling från att enbart vara ett instrument för intern omfördelning till att bli en möjlighet att nylansera och värdesätta relationerna med grannländerna .
herr talman ! från i år står runt 200 miljarder euro till förfogande för strukturfonden fram till år 2006 , men bara 5 3 / 4 procent har reserverats för gemenskapsinitiativen : interreg , leader , urban och equal .
det är en minskning med 3 3 / 4 procent mot hittillsvarande gemenskapsinitiativ .
för equal har inte mer än 2,8 miljarder euro avsatts , vilket framgår tydligt av kollegan ursula stenzels välbalanserade betänkande .
desto mer förvånande är det stora antalet ändringsförslag och den långa önskelistan som rör möjliga uppgifter .
hur skall man då prioritera ?
det råder enighet om grundsatsen att diskriminering och ojämlikheter på arbetsmarknaden skall arbetas bort .
transnationella strategier skall ge eftersatta grupper tillgång till sysselsättning .
jag har ingen förståelse för förslag som innebär att man vill satsa på byråer för utbyte av information om tekniskt bistånd .
dessa byråer var faktiskt föremål för den mest häftiga och berättigade kritik mot den förra kommissionens arbete .
vårt utskott för sysselsättning och socialfrågor gick nu en gång i spetsen för analysen av väsentliga brister och försummelser i kontrollen av leonardo .
kommissionen kan således inte heller när det gäller equal slippa undan det direkta ansvaret och kontrollen . förslag från medlemsstaterna kan kommissionen godkänna endast om dessa uppfyller alla villkor .
för det första : integreringsarbetet genom sektoriella och geografiska utvecklingspartnerskap , varvid hänsyn skall tas till sysselsättningspolitiska grundprinciper . för det andra : systematisk integrering av berörda aktörer , de lokala , regionala och nationella myndigheterna , utbildningscentren , universiteten , de frivilliga organisationerna , arbetsmarknadens parter och den privata sektorn med ett bestående partnerskap som mål .
kommissionen måste alltså förpliktas vad gäller den strategiska ramen för att främja arbetsförmåga och arbetskvalitet , utvärdering av resultaten och den effektiva kommunikationen kring best practices .
först då kan man uppnå den önskade multiplikatoreffekten .
herr talman ! jag vill hänvisa till kommissionens förslag om budgetposten för främjande av den gemensamma jordbrukspolitiken .
den 26 oktober 1999 antog europeiska kommissionen ett förslag för att se till att budgetposten för information till allmänheten om den gemensamma jordbrukspolitiken ( gjp ) får en rättslig grund .
genom detta förslag kommer den befintliga budgetposten b2-5122 att tas bort och en ny budgetrubrik , b1-382 , kommer att skapas .
åtgärder som främjar en förståelse mellan unga jordbrukare och eu , och som också skapar starkare förbindelser med ansökarländerna och resten av världen är viktiga .
jag lägger därför fram dessa ändringsförslag i parlamentet för att detta skall ge sitt stöd till de bidrag som denna typ av program ger .
med beaktande av behovet av att uppmuntra unga jordbrukare att fortsätta driva sin verksamhet , är det oerhört viktigt att de håller sig väl informerade om utvecklingen inom den gemensamma jordbrukspolitiken .
information till och fortbildning av unga jordbrukare på gemenskapsnivå är oerhört viktigt .
jag ber er att stödja att en del av den tillgängliga budgeten skall koncentreras på kunskapsutveckling bland gemenskapens unga jordbrukare .
vad gäller information och fortbildning , så har denna budgetpost tidigare använts för tilldelning av medel till information , kommunikation och fortbildning .
men kommissionen föreslår nu att fortbildning inte längre skall ingå .
jag anser att fortbildning bör ingå i de fall denna ger relevant information om gjp på gemenskapsnivå .
en sådan fortbildning på gemenskapsnivå är ett sätt att se till att unga jordbrukare har den information om gjp som är nödvändig för att kunna fatta bra affärsbeslut för framtiden .
jag lägger därför fram tre ändringsförslag .
jag uppmanar parlamentet att stödja dessa .
jag tar till orda för att , med erfarenhet från den kommunala förvaltningen , uttrycka nyttan av , jag vågar säga nödvändigheten , att urban-programmen har tre inriktningar . för det första att främja återställande av historiska , gamla , kanske ödelagda infrastrukturer och stadsdelar .
för det andra att främja och stimulera den ekonomiska aktiviteten och det sociala livet i dessa historiska kvarter , i dessa delar av de gamla städerna .
vi har ingen större nytta av gator , som nu kanske har utmärkt belysning , med nya trottoarer , med stenbeläggning , kanske vitkalkade och vackra , om vi inte har förmåga att fylla dem med aktivitet och således också sysselsättning .
jag vill förtydliga att det inte handlar om finansiering eller hjälp till olika sociala aktörer utan att också finna en inriktning mot sysselsättning i urvalet av stödberättigade projekt eller , vilket är detsamma , projekt som leder till att gynna skapande av , impulser till och initiativ för sysselsättning .
för det tredje - och kanske skulle man behöva säga att det är det första - , att projektens huvudinriktning måste vara ett fullständigt återvinnande av personer och familjer , eftersom människan inte är gjord för rätten , utan rätten för människan .
i dessa områden i våra städer lever ofta ensamstående föräldrar , äldre som lever på pension och inte längre deltar i produktionen och familjer med svårigheter , ibland upplösta och ostrukturerade .
de bor i områden som borde kunna dra nytta av dessa projekt .
om vi kan uppnå detta med dessa tre inriktningar tror jag att dessa familjer , dessa personer , dessa europeiska medborgare kommer att tro mer på europa och det tycker jag är mycket viktigt eftersom det i slutänden är städerna som kommer att bli mer och mer huvudrollsinnehavarna i det europeiska samhällslivet .
damer och herrar ledamöter ! det är ett egendomligt sammanträffande att vi i dag diskuterar equal-initiativet här i europaparlamentet .
i europa har det den senaste tiden , på grund av den politiska utvecklingen i österrike , funnits en stigande , en ökande politisk oro , det har gjorts politiska uttalanden och förekommit politiskt samtal .
det bör betonas att såväl parlamentet som kommissionen har lagt fram särskilda strategier .
särskilda förslag såväl om lagstiftning som om åtgärdsprogram som avser bekämpningen av diskriminering , som avser uppbyggnaden av samhällen med friheter och lagar .
så , jag nämner helt kort paketet mot diskriminering och ber med anledning av det att de respektive ansvariga parlamentsutskotten utser föredragandena , så att vi så snabbt som möjligt kan gå vidare med paketet mot diskriminering .
och jag kommer till equal-initiativet , som naturligtvis grundar sig på artikel 13 .
equal-initiativet avser alla former av diskriminering på grundval av artikel 13 , det vill säga bekämpning av diskriminering som grundar sig på ras , kön , ålder , handikapp .
jag skulle särskilt vilja tacka stenzel , för hennes arbete med att försöka nå en överenskommelse om equal-initiativet är enastående svårt och komplicerat , såväl på grund av att utskott som ser på saken ur en annan synvinkel är inblandade som på grund av att det är en enastående känslig politisk fråga .
min första kommentar , som även har formulerats av många kolleger , gäller frågan om huruvida kvinnorna måste tas upp separat .
jag håller med om att det i artikel 13 finns en sak som vi inte håller med om , men fördraget är sådant i dag , och bland diskrimineringskategorierna finns på lika bas även diskriminering som grundar sig på kön .
med fördraget som grund , i den form som det har i dag , är equal-initiativet sammansatt på det sättet .
jag vill dock påminna om att det finns en särskild pelare i sysselsättningsstrategin som gäller kvinnorna och att ett särskilt program , det femte programmet för jämlikhet mellan män och kvinnor , håller på att förberedas .
jag har indelat frågorna som damerna och herrarna parlamentskolleger har berört i fyra grupper
för det första , utvidgningen av de tematiska enheterna .
det finns fyra tematiska enheter , liksom i sysselsättningsstrategin : anställbarhet , företagaranda , anpassningsförmåga och lika möjligheter , och vi instämmer i utvidgningen av dessa tematiska enheter i enlighet med de förslag som har lagts fram av europaparlamentet .
angående oron över risken att ett land lägger alla pengar på en av de kategorier som är utsatt för diskriminering , skall jag säga att det klart och tydligt sägs i initiativet att medlemsstaterna bör presentera en tematisk kategori för var och en av de grupper som är utsatta för diskriminering .
den andra frågan gäller flexibilitet och förenkling .
jag håller med leinen om att språket i initiativet verkligen är mycket svårt och ogenomträngligt .
av den anledningen håller avdelningarna redan nu på att revidera texten , att förenkla dess struktur och göra dess språk mer lättförståeligt .
angående frågan om flexibilitet , vill vi med vårt förslag få till stånd utvecklingspartnerskap och utvecklingssamarbete , såväl på geografisk nivå , där grupper av olika slag skall samarbeta i en bestämd geografisk region för att bemöta diskriminering på arbetsområdet , som på tematisk nivå , där det till exempel skall kunna förekomma samarbete i en konkret ekonomisk sektor .
här kommer det att finnas ett stort utrymme för flexibilitet i medlemsstaterna , och de kommer att kunna anpassa utvecklingssamarbetet i enlighet med sina önskemål .
en förutsättning är naturligtvis att medlemsstaterna samarbetar och att vi har ett nät med vars hjälp vi kan utbyta erfarenheter .
avslutningsvis skall jag ta upp det tekniska biståndet .
vi vill att det skall finnas fyra stödkategorier .
för det första skall förberedelserna stödjas , för det andra genomförandet , för det tredje samarbetet mellan aktörerna , så att ett erfarenhetsutbyte kommer till stånd , och för det fjärde det tekniska biståndet .
eftersom det har funnits ett stort engagemang och en stor oro över frågan om hur det tekniska biståndet skall tillhandahållas , skall vi säga att externa byråer kommer att användas .
det är omöjligt , vilket också min kollega barnier sade , att kommissionens tjänstemän skall utföra allt det arbete som fram till i dag har utförts av externa medarbetare .
målet är att det på nationell och europeisk nivå skall finnas stora grupper av åtgärder som offentliggörs , och det kommer att finnas en fullständig beskrivning av det arbete för vilket det externa biståndet begärs och en fullständig beskrivning av den produkt som vi förväntar oss av varje teknisk byrå , så att det är möjligt att både övervaka och utvärdera detta arbete .
jag vill understryka att det är enastående viktigt att det aktuella initiativet främjas så snabbt som möjligt , dels på grund av politiska omständigheter , men även på grund av att vi anser att det är viktigt att det träder i kraft som planerat , dvs. att vi måste vara helt förberedda i slutet av 2000 .
justering av protokollen från de två föregående sammanträdena
protokollen från sammanträdena torsdagen den 3 februari och måndagen den 14 februari har delats ut .
protokollet från den 3 februari delades i själva verket ut redan i bryssel . det är kanske därför som en del kolleger inte hade fått det .
( prokollet justerades . )
tack , herr medina ortega .
jag delar fullt ut det beklagande som ni uttrycker .
skulle ni vänligen vilja skriva till mig så att jag med stöd av bevis kan anmäla detta till de behöriga ansvariga såväl hos air france som den franska regeringen ?
jag tror verkligen att det inte längre är möjligt och att vi absolut måste protestera med full energi .
fru talman ! igår upplevde jag och medina ortega samma sak .
jag tycker att de franska myndigheterna - som har äran att hysa europaparlamentets säte i strasbourg - bör vara medvetna om sitt ansvar för att garantera fungerande kommunikationer med alla unionens huvudstäder .
just det , herr napolitano , tack för det .
fru talman ! det handlar här inte om försenade plan : jag skulle vilja be om ursäkt för min kollega i gruppen de gröna , caroline lucas , som är brittisk ledamot .
hon kunde inte närvara eftersom hon hade arresterats vid en demonstration mot kärnkraft i glasgow i går morse .
hennes identitet noterades : det framkom mycket tydligt att hon är ledamot av europaparlamentet , ändå kvarhölls hon i arrest hela dagen .
jag anser att det är absolut oacceptabelt och jag ber er - jag har för övrigt skrivit till er tillsammans med min kollega hautala i det avseendet - intervenera hos de brittiska myndigheterna för att sådana händelser inte skall upprepas och att man ber lucas om ursäkt .
tack , herr lannoye .
jag har fått er skrivelse och har redan vänt mig till den brittiska delegationen .
fru talman ! med tanke på omröstningen i dag vill jag be om något som jag berörde redan i går vid debatten om equal-betänkandet .
jag ber om att man uppskjuter omröstningen i dag om gemenskapsinitiativet equal , eftersom vi helt enkelt behöver litet mer tid för att komma överens om en viktig punkt .
jag är optimistisk och ser verkligen med lugn och tillförsikt fram emot omröstningen ; vi kommer att få ett synnerligen brett godkännande av detta yttrande om equal .
vi behöver bara litet mer tid för att utarbeta detaljerna i samband med asylfrågan , och jag ber därför om att omröstningen genomförs i morgon i stället för i dag .
fru talman ! för att fortsätta från den punkt som lannoye tog upp : lucas arresterades precis utanför glasgow för att hon protesterade mot tridentbasen i faslane .
jag sympatiserar mycket med den protesten .
jag har dock ingen sympati för lucas som försöker gömma sig bakom sin parlamentariska immunitet .
jag har också varit arresterad för att ha protesterat i faslane .
jag gömde mig inte bakom någon immunitet .
jag tog det straff som jag fick .
lucas borde göra detsamma .
fru talman ! jag skulle vilja kommentera stenzels yrkande om att skjuta upp omröstningen om gemenskapsinitiativet equal till i morgon .
detta initiativ har faktiskt diskuterats mycket livligt i utskottet , och eftersom det är ett viktigt förslag från kommissionen , som gäller de överenskommelser vi träffade förra året , tycker jag att det kan antas .
vi är överens med stenzel om att yrkandet om uppskjutande kan bifallas för att finna största möjliga samförstånd mellan grupperna , så att parlamentet med bredast möjliga majoritet uttrycker sin ståndpunkt om detta initiativ .
finns det några kolleger som vill yttra sig mot stenzels begäran , som ghilardotti just stödde ?
eftersom det inte är så , tar vi upp den till omröstning .
fru talman ! enligt artikel 29.4 skall ni hållas informerad av de politiska grupperna om varje ledamot som anslutit sig till en ny politisk grupp eller lämnat en politisk grupp .
har ni fått någon anmälan om att några medlemmar lämnat gruppen europeiska folkpartiet eller tillhör österrikiska folkpartiet fortfarande denna politiska grupp ?
herr corbett , jag har inte hört talas om någonting .
när det gäller föredragningslistan för torsdagen föreslår jag er , mot bakgrund av en begäran som inlämnades i går vid plenarsammanträdet , att förlänga debatten om brådskande och aktuella frågor med en halvtimme , det vill säga fortsätta fram till kl. 18.00 . omröstningen kommer att äga rum kl. 18.00 .
strategiska mål och lagstiftningsprogram från kommissionen
nästa punkt på föredragningslistan är den gemensamma diskussionen om kommissionens uttalanden om sina strategiska mål för en femårsperiod och om det årliga lagstiftningsprogram för år 2000 .
fru talman , ledamöter ! ett femårsprogram är ett viktigt åtagande och därför tyckte jag det var bättre att ni alla fick hela texten till talet utdelad , den finns på fyra språk .
för att respektera tidsbegränsningen skall jag endast ta upp de stora dragen i mitt program : ett program för början av en mandatperiod och för början av ett nytt sekel under vilket man har både rättighet och skyldighet att se europa i ett vidare perspektiv , ett europa som för närvarande upplever en motsägelsefull tid .
vi skall komma ihåg att europa under sina femtio års historia har gett oss fred , säkerhet och frihet , och att det enade europa också har bidragit till att ge oss en period med aldrig tidigare skådat välstånd .
nu känner vi av början på en solid återhämtning som även verkar kunna bli mycket varaktig om vi för en klok politik , en återhämtning som är en logisk följd av de ansträngningar vi har gjort .
vi får den inte gratis , utan som en konsekvens av saneringen av de offentliga finanserna i europas länder , som har hållit inflationen under kontroll med en klok politik inriktad på kostnadskontroll och ökad produktivitet . detta i ett europa som har inlett en energisk omstrukturering av sina industrier , banker och sin offentliga service , även om denna process ännu inte är fullbordad , även om det fortfarande är långt kvar att gå .
trots dessa aspekter finns det ändå besvikelse och oro i europa : besvikelse och oro för arbetslösheten som inte minskar tillräckligt snabbt , för en teknisk eftersläpning som framstår som större och större , och som framför allt börjar åtföljas av en kraftig eftersläpning också inom det vetenskapliga området , för de europeiska institutionerna som verkar vara långt efter , som inte verkar vara tiden vuxna , i första ledet kommissionen själv .
kommissionen kris var faktiskt en avgörande punkt i förhållandet mellan europa och dess medborgare , och det låga valdeltagandet i europavalen var ett oroande tecken på detta .
något som går ännu djupare är dock känslan av osäkerhet , känslan av att inte vara förberedd för den nya värld som växer fram , en värld som förändras totalt , som genom globaliseringen kommer att förändra också våra referensramar .
detta är ingenting alldeles nytt i historien : europa har redan tidigare en gång genomgått en liknande förändring med en explosionsartad ökning av marknaderna , förändrade referensramar och en ny världsuppfattning .
jag syftar på femtonhundratalet , efter upptäckten av amerika , då allting förändrades .
vissa länder - såsom frankrike och spanien - visste att svara på utmaningen och gav upphov till stora nationalstater . andra länder - såsom italien - klarade inte denna utmaning och förlorade all den dominans de hade byggt upp under millenniets första hälft : en dominans inom vetenskap , teknologi , ekonomisk utveckling , försvarsstrukturer och militär organisation , filosofi och litteratur .
i dag står europa inför en liknande utmaning och vi vet att historien kommer att vara lika skoningslös som förr i tiden .
mot bakgrund av dessa stora förändringar fordras ett ekonomiskt starkt europa för att förhindra att våra nationalstater även nu försvinner genom en globalisering med dimensioner och utmaningar utan motstycke i vår historia . globaliseringen påbjuder nämligen enhet .
varje dag hör vi nyheter om nya avtal på global nivå och varje dag hör vi nyheter om förändringar också på europeisk nivå . men ännu mer nödvändigt är att europa känner sig starkt på det politiska planet .
tidigare har den inre marknaden och den gemensamma valutan varit den fasta punkten i vårt handlande , det bärande elementet i europas liv .
i dag är de nya gränserna för den europeiska integrationen politiska gränser : den gemensamma utrikes- och säkerhetspolitiken , den inre rättvisan och säkerheten och - på ett underordnat plan - den avgörande frågan om de grundläggande politiska värderingar vår samexistens vilar på .
därför har kommissionen antagit den strategiska planen för 2000-2005 , en plan som genast översändes till europaparlamentet , som ni redan känner till och som jag alltså inte skall beskriva i detalj här .
någon kanske anser att den är för allmänt hållen , men inga politiska instanser upprättar detaljerade femårsplaner .
detta är europeiska unionen , inte sovjetunionen .
i vår plan anges de stora referensramarna , vår verksamhets inriktning i stort : för det första att utveckla nya styrelseformer för europa , för det andra att expandera och utvidga området för fred , frihet och säkerhet , för det tredje att lansera en ny ekonomisk utvecklingsfas , för det tredje att värna och öka livskvaliteten .
dessa är våra stora handlingslinjer för de kommande fem åren .
vad den första beträffar - de nya styrelseformerna för europa - vet ni redan att kommissionen har åtagit sig att lägga fram en vitbok och inte en komplett lagtext eftersom kommissionen inför de stora frågor som förändrar strukturen för vårt umgänge först tar fram ett debattunderlag . sedan diskuterar vi innehållet med er , och ur detta uppstår ett först politiskt dokument och slutligen en lagtext .
detta är ett öppet och kraftfullt sätt att gå till väga , så att alla europeiska institutioner och europas befolkning involveras .
denna vitbok är ett svar på de utmaningar utvidgningen ställer upp . det är utvidgningen som tvingar oss att se över hur alla våra institutioner fungerar , att till och med se över vår politik - all vår politik - och framför allt tänka igenom vad vi skall fortsätta att göra på unionsnivå när medlemsländerna är tjugofem eller trettio , vad som bättre görs av de enskilda staterna , regionerna eller de lokala myndigheterna .
men det är inte bara utvidgningen som driver oss till denna översyn : som jag sade nyss är det också globaliseringen av ekonomin och politiken .
vi måste styra europa så att vi blir mer effektiva , kommer närmare medborgarna och verkar för allas delaktighet . först och främst måste vi ta itu med den stora frågan om kvinnors delaktighet .
i den jämförelse mellan europa och förenta staterna som nyligen gjordes är en av de stora skillnaderna inte så mycket arbetskraftens rörlighet eller tillgången på riskkapital utan kvinnors deltagande i det ekonomiska livet , ett deltagande som i förenta staterna har helt andra dimensioner än i europa .
det handlar om ett område där europa tvärtom alltid har varit ledande : detta måste vi alltså tänka igenom på djupet och öppet , och alla institutionerna - kommissionen , parlamentet och rådet - måste tänka igenom sin roll och sin politik .
vi kommer alltså att omedelbart börja arbeta med denna vitbok , även om vi måste avvakta resultaten fån regeringskonferensen innan vi slutför den och den därför inte kan läggas fram förrän våren 2001 .
det blir ingen filosofibok utan en konkret bok med många detaljerade förslag .
vi - kommissionen - är de första att veta att vi måste göra en total översyn av oss själva , och därför kommer vi att göra två saker : vi kommer att engagera oss och vi engagerar oss redan nu till fullo i den interna reformen , och vi kommer att tänka igenom vår politik på djupet .
jag har bett alla kommissionärer - och vi kommer att be dem om en ännu djupare analys - att identifiera all verksamhet som kan läggas ned .
kommissionen måste fastställa sin kärnverksamhet , den verksamhet vi skall koncentrera oss på , och upphöra med mindre viktig verksamhet för att frigöra nya resurser och få ett korrektare och mer samarbetsbetonat förhållande med de enskilda länderna , med regionerna och med de lokala samhällena .
vi skall alltså frigöra nya resurser , men det kommer också en tid - fruktar jag , och jag vill säga det här inför parlamentet - då även dessa nya resurser som vi redan håller på att frigöra inte kommer att vara tillräckliga för att vi skall kunna ta itu med våra nya uppgifter : jag tänker på utvidgningen , på den nya rättsliga och inrikespolitiska sektorn , på hälso- och sjukvårdsfrågorna , på miljöfrågorna .
den dagen , när vi har utnyttjat alla våra resurser maximalt , kommer jag inte att tveka att inställa mig inför er för att be om nya resurser , men jag säger redan nu att om vi inte har erforderliga resurser måste vi vägra ta på oss några nya uppgifter , eftersom det inte finns någon överensstämmelse mellan de nya uppgifter vi tar på oss och de resurser vi har till vårt förfogande .
vad den interna reformen beträffar känner ni väl till det engagemang min kommission har lagt ned på denna fråga från första dagen .
jag vet mycket väl att vi inte kan uppnå några politiska mål om kommissionen inte reformerar sig internt kraftigt och genomgripande , om vi inte blir effektivare , om vi inte tar ett effektivitetssprång inom alla sektorer med början i den sektor där vi hittills har samlat på oss den mest dramatiska eftersläpningen , det vill säga inom det externa biståndet .
att ge hjälp snabbt när den behövs räddar människoliv . att ge den för sent kan i många fall vara värre än att inte ge den alls .
när jag talar om externt bistånd går mina tankar i första hand till balkan , där det finns en stråle av hopp tack vare våra funktionärers engagemang på fältet , ett extraordinärt engagemang med tanke på de organisatoriska problem vi har .
jag tänker även på bernard kouchners bemödanden , på stabilitetspakten som vi står bakom med kraft , med total hängivelse , men jag tänker också på de nya händelserna i till exempel kroatien , där situationen har förändrats på några veckor : de europeiska institutionerna öppnade omedelbart dörren för en dialog med detta land , de mottog denna nyhet väl medvetna om att inte bara bosniens utan framför allt serbiens problem endast kommer att kunna lösas om vi slår en demokratisk järnring kring serbien .
detta är det nya element vi måste bidra till att införa på balkan .
vi måste bli effektivare på detta område , vi måste öppna donau för trafik igen .
det är motsägelsefullt att erbjuda hjälp till rumänien och bulgarien och låta dessa länders stora resurs vara blockerad .
vi måste rena floden och därför kommer den miljöansvariga kommissionären under de närmaste dagarna att lägga fram detaljerade projekt för att få bukt med detta allvarliga problem .
vi har gjort mycket på balkan : den nya europeiska byrån för återuppbyggnad av kosovo , insatsstyrkan för balkan , en ny förordning för att snabba upp rutinerna . vi måste dock absolut göra mer .
vi måste liberalisera handelsutbytet inom regionen och utbytet mellan denna region och europeiska unionen .
vi måste bidra till att konstruera infrastruktur som bryter en sekellång isolering . vi måste intensifiera ansträngningarna för att i dessa länder bygga upp demokratiska och pluralistiska samhällen med ett civiliserat samhälles institutioner , offentliga strukturer , ordningsmakt och organisation , men framför allt måste vi få dessa länder att arbeta tillsammans och se regionen som en enhet både politiskt och ekonomiskt .
om vi inte gör det har vi misslyckats med vår uppgift .
minns att marshallplanen på sin tid inte bara hade effekt på grund av sina stora resurser : den fick ännu större effekt eftersom den tvingade oss européer att arbeta tillsammans med ett nytt perspektiv , att ge vår politik och vår ekonomi en ny horisont .
detta är vad vi måste göra för balkan .
europa måste för balkanländerna och hela resten av världen bevisa sin förmåga att utvidga området för säkerhet , fred och frihet , sin kapacitet att spela en huvudroll på den internationella scenen .
självfallet kommer vi åter igen tillbaka till utvidgningen , som måste genomföras genom att man samtidigt utvidgar området för säkerhet , fred och frihet .
vi har lovat mycket i denna riktning men jag tror att vi kommer att kunna hålla våra löften även om vi har en mycket delikat uppgift framför oss .
utvidgningen , som kommer att följa oss under hela vår femårsperiod och även senare - jag tänker på kandidatländernas förhoppningar - måste komma till stånd med säkerhet och objektiva kriterier , men den måste också komma till stånd så att man lugnar den allmänna opinionen i de berörda länderna och , än mer , lugnar vår egen allmänna opinion .
det kommer att bli vänskap , harmoni och öppenhet , men också stränghet i utvidgningen .
jag upprepar : vi måste lugna den allmänna opinionen i de länder som vill bli medlemmar , men vi måste lugna vår egen allmänna opinion ännu mer .
våra skyldigheter upphör inte med utvidgningen , de upphör inte med balkan .
det finns några andra frågor som är avgörande : förhållandet med ukraina , förhållandet med ryssland , förhållandet med våra grannländer och i än högre grad den stora frågan om förhållandet med södra medelhavsområdet , som kommer att bli den avgörande punkten i den europeiska historien , för kommande generationers säkerhet och trygghet i europa .
i denna mening har vi en skyldighet mot hela afrika : afrika som man har vänt sig till med förhoppningar på den senaste tiden , som har fått mottaga erbjudanden men där ännu ingenting konkret har genomförts .
afrika där övergången under de senaste åren inte har varit från totalitära regimer till demokrati utan tvärtom , från demokrati till totalitära regimer .
afrika som är bekymmersamt för oss att konfronteras med .
därför har vi ytterligare en uppgift på det internationella planet , vilken kommissionären med ansvar för handelsfrågor redan har föreslagit : uppgiften att återuppta millennium round , med ett stort tillmötesgående som vi redan tagit på oss och erbjöd redan innan seattle , men som inte kunde konkretiseras . att alltså ta över bördan för vissa grundläggande problem från de fattigaste länderna , inte bara vad gäller avskrivning av skulder utan även att ensidigt öppna för handel med världens fattigaste länder .
det krävs en ny lösning , annars kommer händelser som de i seattle alltid att upprepas och förhindra att europa utövar en positiv roll i historien .
överallt i världen måste europas agerande styras av stor respekt för principerna om frihet , respekt för individens rättigheter och respekt för minoriteters rättigheter .
låt oss komma ihåg att vi , europeiska unionen , är en union av minoriteter : alla vi är i minoritet i europa .
det finns en oro även hos våra femton länder , en oro som kanske kommer att uppstå igen under den kommande tioårsperioden .
jag talar om fallet österrike , där kommissionen har varit sin roll trogen . vi har verkat för sammanhållning av unionen men varit orubbliga i vårt försvar av fördragen , redo att bestraffa varenda litet övertramp som innebär ett brott mot principerna om demokrati , rättigheter och respekt för minoriteter .
vissa har kritiserat mig för det lyckönskningsmeddelande jag skickade till kansler schüssel .
jag skall säga er : förväxla inte en nödvändig och pliktskyldig formell hövlighet med mindre reell fasthet .
läs brevet igen : hänvisningen till unionens grundläggande värderingar är ett utdrag ur fördragets artikel 6 , jag upprepar artikel 6 i fördraget , och detta är ingen tillfällighet .
jag frågar er också : tror ni att kommissionen någonsin har påmint någon annan nyvald europeisk regeringschef om dessa principer ?
det är detta vi vill göra : bibehålla vår roll av övernationell struktur , bibehålla den roll vi har fått genom fördragen , men också vara obevekliga om principerna och utgå från fakta i våra bedömningar .
i november förra året lade kommissionen fram ett förslag till direktiv mot rasismen .
jag ber rådet att snabbt anta det och jag ber parlamentet att hjälpa oss i denna kamp , som ytterligare fördjupar den grundläggande basen för vår sociala sammanhållning .
jag skall avsluta med att snabbt påminna om de sista två punkterna i vårt program : ekonomin och livskvaliteten .
jag har redan talat om ekonomin : vi är väl medvetna om vilka grundingredienserna är för att föra in europa på vägen mot en återhämtning som kan vara länge och äntligen skapa arbetstillfällen .
vi måste fortfarande hålla inflationen nere , fortsätta med avregleringen , värna konkurrensen i än högre grad , driva på spridningen av informationsteknologi och av all ny teknik , driva på vetenskapen , vetenskapens förfront , njuta av att befinna oss i vetenskapens förfront .
det kommande toppmötet i lissabon om dessa frågor - spridning av teknik och sysselsättningen - blir ett avgörande toppmöte .
det behövdes fyra år innan vi kunde ha ett toppmöte av detta slag .
nu kommer vi äntligen att ha det : vi får inte missa tillfället .
det sista åtagandet är slutligen att öka livskvaliteten .
vi inledde detta kapitel med vitboken om livsmedelssäkerhet : nu måste vi göra stora framsteg på miljöområdet .
fallet med fartyget erika och giftutsläppet i donau visar hur angeläget det är med insatser på europeisk nivå till skydd för miljön .
det är dags att fundera på , och sedan förverkliga , en europeisk räddningstjänst .
i allt för många fall hör man krav på detta efter det att katastrofen har inträffat .
jag tror att man måste börja tänka på dessa saker innan katastroferna inträffar .
dessa är de utmaningar vi har framför oss : vi som kommission men också alla de andra europeiska institutionerna .
ledamöter , fru talman , hur skall vi mäta våra fem verksamhetsår ?
hur skall vi mäta resultaten av dessa fem år ?
jag vet inte , men en måttenhet kan helt klart vara den kamp vi måste utkämpa tillsammans .
låt oss ta en mycket enkel parameter : valdeltagandet vid nästa europaval .
om det blir högre än vid det föregående valet betyder det att vi har vunnit vår kamp .
fru talman , ärade ledamöter ! vi har alla dessa stora politiska utmaningar framför oss , men vi har också stora möjligheter framför oss , just på grund av den återhämtning som har inletts .
detta , ärade ledamöter , kan bli europas decennium .
jag säger : detta måste bli europas decennium .
fru talman , herr kommissionsordförande ! jag vill börja med att välkomna denna framställning av och unika debatt om regeringens - ett ord som ordförande prodi och även jag är förtjusta i- kommissionens program för hela mandatperioden .
i första hand för att det innebär att vi kan förklara för våra medborgare vad vi har för avsikt att göra och vad vi redan håller på att göra .
dessutom måste vi beklaga och med tanke på framtiden försöka rätta till den nuvarande situationen : det har tagit oss nästan elva månader - ordförande prodi blev föreslagen på toppmötet i berlin i mars i fjol - att skapa ett lagstiftningsprogram .
felet är inte enbart hans ; vi håller på att övervinna en kris , men jag anser att det lämpligaste , med tanke på framtiden , är att tillsättandet av nästa kommission sammanfaller med framläggandet av ett lagstiftningsprogram .
vi håller på att göra förändringar , men situationen är komplicerad .
ordförande prodi inledde sitt tal genom att ta upp en paradoxal situation , en paradox inom europeiska unionen och även i världen som sådan : vi står på tröskeln till ett nytt konfessionslöst årtusende , som styrs av spindelnätet internet och de biotekniska framgångarnas häxkonst ; faktum är att vi upplever övergången till en ny epok , men om vi begränsar oss till det som i dag är europeiska unionen och talar om regeringar och regerande - som åtminstone på spanska för tankarna till det tidigare namnet på inrikesministeriet , men kanske är det också intressant att tala om regerande - , så är det viktigaste att europeiska unionen får en bra regering och eftersom ordförande prodi alltid försvarar sin födelseort bologna , råder jag honom att åka till siena för att ta sig en titt på något som vi alla begriper oss på , nämligen ambrogio lorenzettis fresker , där han skildrar bon governo och mal governo .
det vi behöver här är en bra regering , fru talman .
eftersom vi håller på att hämta oss efter en mycket svår kris , måste vi försöka fylla våra institutioner med innehåll och lyfta fram dessa .
jag vill för parlamentet nämna ett faktum som vi ofta glömmer , nämligen att tillsättandet av prodis kommission i september förra året vann starkt stöd i omröstningen , något som enligt vår uppfattning är tecken på en reformvänlig och europavänlig majoritet .
jag vill emellertid påpeka att man i samband med denna breda överenskommelse i vissa grupper sade att majoriteten av parlamentet bör utgöra en opposition till en majoritet i rådet .
det skulle utgöra ett hinder för något viktigt , nämligen utvecklandet av medbeslutandet i lagstiftningsprogrammet .
jag påpekar detta , eftersom jag anser att stödet till kommissionen måste ske kontinuerligt under hela mandatperioden .
å andra sidan får vi ta del av det politiska europas födelse , en gemenskap med värderingar som vi delar , en europeisk union i medborgarnas tjänst .
vad beträffar den senaste tidens händelser vill jag säga - och det kommer jag att säga den dag eller i början av den vecka som regeringskonferensen inleds - att vi verkligen måste lägga större vikt vid och lyfta fram arbetet med stadgan för de grundläggande rättigheterna som jag , efter det som vi har sagt till följd av den österrikiska krisen , absolut anser bör ingå i fördragen .
jag tvivlar inte ett ögonblick på detta och ser det som en viktig faktor .
därför , fru talman , vill jag även påpeka att vi måste vara medvetna om och försiktiga med vårt språkbruk .
förra veckan beskrev den österrikiska koalitionens nya finansminister det österrikiska parlamentet som en komedi och en teater .
vi som har tvingats leva under en diktatur vet att en diktatur kan råda med ett skuggparlament .
däremot är det ingen demokrati utan ett levande parlament .
jag tror att ett sådant språkbruk är extremt farligt , och fördömer härmed detta .
vad beträffar de fyra viktigaste prioriteringar som ordförande prodi ständigt hänvisar till , vad beträffar analysen av de utmaningar som väntar , vill jag påstå att vi är helt överens .
jag vill ändå påpeka för kommissionen att den socialistiska gruppen har förändrat sin syn på prioriteringarna .
vi uppfattar det som att den första prioriteringen är den ekonomiska och sociala agendan , som inbegriper det som i era prioriteringar kallas livskvalitet , det vill säga medborgarnas rättigheter som konsumenter och även som individer i förhållande till sådant som vi alltid bekräftar , men som vi inte poängterar tillräckligt , så som den europeiska sociala modellen och anpassningen av den till nya situationer , konsumenternas rättigheter samt respekten för miljön och en hållbar utveckling .
när man talar om löftet om full sysselsättning , måste utgångspunkten vara att full sysselsättning i dag inte , som på beveridges tid i slutet av andra världskriget , enbart innebär sysselsättning för familjens manliga överhuvud .
vi måste bekräfta jämlikheten mellan könen , den så omtalade gender mainstreaming , som är en av de punkter som är minst utvecklad i kommission prodis program .
det förutsätter en prioritering av jämlikheten mellan könen , en anpassning av den sociala modellen och i synnerhet en tydlig kamp mot populismen i ett läge då vår ekonomiska och sociala sammanhållning är hotad , och det bör också vara den främsta prioriteringen i kommissionens arbete .
det bör förstärkas genom en tydlig kamp mot rasism och intolerans , så att man i praktiken bekräftar framväxten av en union som numera har en stark attraktionskraft på den övriga världen och som har förvandlats till ett område för immigration tack vare sin framgång och befolkningens höga medelålder .
jag anser att det är det första mål vi bör uppnå .
i det sammanhanget vill jag nämna ytterligare en faktor , nämligen den ekonomiska regeringen med en gemensam valuta - jag tror att den kommer att slå igenom- och även på den punkten måste kommissionen göra framsteg .
jag skulle vilja ha - det vill säga min grupp skulle vilja ha - en större tydlighet vad beträffar granskningen av agenda 2000 , angående de ambitiösa målsättningarna och i synnerhet något så viktigt som kommissionen har gjort , nämligen att anamma utvidgningen i förhandlings- och integrationsprocessen .
föreställer sig kommissionen en granskning först i slutändan ?
frågan om beskattning betraktar vi också som en nyckelfråga .
vad gäller regerandet i allmänhet , kan det vara intressant att göra vissa teoretiska överväganden .
en sak vill jag påpeka : det är farligt att härifrån ompröva europeiska unionens regerande .
jag är definitivt en anhängare av subsidiaritetsprincipen .
om vi lyckas definiera det område vi skall regera inom , tror jag att det skulle vara mycket positivt .
för övrigt anser jag att våra överväganden även skall gälla subsidiaritetsprincipen .
detta ska inte enbart gälla kommissionen - även våra stater , våra parlament och vårt civila samhälle måste överväga subsidiaritetsprincipen .
slutligen , fru talman , vill jag kort hänvisa till det sista mål , som enligt vår uppfattning är högst grundläggande : en stabilisering av kontinenten och ett stärkande av europas roll i världen .
på den punkten vill jag påstå att det råder enighet och att det finns ett stöd vad gäller prioriteringen av sydöstra europa , utvidgningen och - det har jag redan påpekat - integrationsprocessen och stärkandet av programmet europa-medelhavsländerna samt av vår förmåga att förebygga konflikter , och en fråga som diskuteras mycket , nämligen utmaningen norr-söder .
vi får inte glömma afrika som är den kontinent som inte bara gud utan även europa glömde , inte heller vårt viktiga bidrag till utvecklingssamarbetet .
och slutligen ett område på vilket vårt ansvarstagande ständigt växer , som världens främsta ekonomiska och kommersiella maktfaktor , nämligen som europeiska unionens röst i världen , något som inte bara förutsätter en aktiv attityd inför millennierundan .
det förutsätter även en reform av förenta nationerna och av de internationella finansinstituten , och där har europa ett enormt ansvar .
framför allt måste vi , fru talman och mina damer och herrar , kunna ge uttryck för detta i tydliga ordalag genom att i vissa avseenden ändra den jargong som vi använder oss av , för vi kan inte förvänta oss att européerna , som lever i en tid av genomgripande förändringar , skall ansluta sig till oss med entusiasm om vi fortsätter med ett internt språkbruk över deras huvuden .
det är den främsta metoden att öka och stärka det förtroende som jag hoppas , i vilket fall som helst kommer att kunna mätas i nästa europaval .
fru talman , ärade kommissionsordförande ! jag värderar högt den öppenhet med vilken ni medger att unionen i grunden måste ändras .
ni dryftar mycket grundläggande frågor i ert program .
jag tror att medborgarna börjar intressera sig mera för politik om vi tar fram stora frågor vid sidan av de små vardagliga ärendena .
samtidigt måste man dock säga att ert program i många avseenden tyvärr påminner om ett partiprogram .
det innehåller nämligen många goda avsikter men saknar i stor utsträckning konkreta förslag på hur allt detta skall genomföras .
liksom vilket partiprogram som helst innehåller det också många inre motsättningar .
jag skulle genom mitt eget inlägg vilja hjälpa er att identifiera dessa inre motsättningar .
för det första angående ekonomin och den sociala utvecklingen : man måste kunna dryfta hur vi skall förena målsättningarna för konkurrens med dem för full sysselsättning ; detta omnämns ju i ert program .
borde man när allt kommer omkring utveckla ett konvergenskriterium där man - vilket ni faktiskt antyder i detta program - ställer upp som mål att arbetslösheten inte i något medlemsland får vara högre än i låt oss säga de tre länder som lyckas bäst i den här saken ? en ekologisk skattereform är det som min grupp vill prioritera .
vi kan nämligen skapa sysselsättning och hållbar utveckling endast genom att ändra skattestrukturen , men tyvärr är detta - som vi alla vet - ett område där europeiska unionen är helt oförmögen att handla .
var vänliga och ta upp denna fråga på regeringskonferensen .
europeiska unionen erhåller befogenheter endast genom att koncentrera sig på uppgifter som de enskilda länderna inte kan sköta på egen hand .
i det här avseendet delar säkert parlamentet er uppfattning om vikten av överstatligt beslutsfattande .
en inre motsättning i ert program berör globaliseringen .
jag tycker det är mycket bra att ni tar upp begreppet &quot; global kontroll &quot; , liksom också andra här har konstaterat .
tag dock även lärdom av händelserna i seattle : man måste förena å ena sidan fri världshandel och å andra sidan allt det ur mänsklig synvinkel värdefulla som vi vill värna om .
ni måste inleda en dialog med medborgarsamhället .
var vänliga och demokratisera de internationella organisationerna .
europeiska unionen skulle kunna spela en avgörande roll i den process , där förenta nationerna och världshandelsorganisationen verkligen ställs under demokratisk kontroll .
vi kan lägga fram motioner om detta tillsammans med er .
slutligen ser jag det som mycket positivt att ni så ofta talar om medborgarsamhället , men detta utgör tyvärr en inre motsättning .
ni borde också dra slutsatser vid regeringskonferensen .
man måste ta initiativ så att medborgarna verkligen direkt kan påverka beslutsfattandet .
det ni nyss sade oss är alldeles sant : människorna vill ha en mera aktiv demokrati .
detta är enligt min mening den enda möjligheten om vi vill att folk skall acceptera europa och intressera sig för europa .
fru talman ! min grupp var bland dem som ville ha ett dokument för att snarare kunna ha ett utbyte inom gruppen om kommissionens strategiska mål före debatten än att bara kunna avge en direktreaktion på ett uttalande i plenarsammanträdet .
den främsta fördelen med texten i detta meddelande är således , enligt vår åsikt , att den finns till .
vi är dessutom inte likgiltiga för vissa påståenden som görs i den eller avsikter som framförs , och som prodi i sin tur just har understrukit och rent av klargjort i vissa punkter på lämpligt sätt .
ja , den aktuella globaliseringsprocessen är , jag citerar &quot; snarare uteslutande än inbegripande och har ökat orättvisorna &quot; och därmed bör europeiska unionens ambition vara att bidra till , jag citerar igen , &quot; att nya spelregler fastställs inom unionen och i de internationella förbindelserna &quot; .
ja , många av våra landsmän är , jag fortsätter att citera , &quot; modlösa och ångestfyllda &quot; , för att de inte får se verkliga och hållbara lösningar på väsentliga eller existentiella problem såsom arbetslöshet och social uteslutning vilket påminner oss om det som bör vara en av våra absoluta prioriteringar .
ja , vi måste tänka om i fråga om många aspekter av den aktuella gemenskapspolitiken om vi vill lyckas med det stora men svåra utvidgningsprojektet och vi behöver också , jag citerar , &quot; ha rent strategiska partnerskap med våra grannar från söder och från öster för att bidra till stabilitet och fred &quot; .
vi saknar då inte områden på vilka vi kan inleda allvarliga diskussioner .
vi kommer att noggrant granska de anmälda vitböckerna och på ett konstruktivt sätt delta i de mångtaliga påbörjade och utlovade uppbyggnadsplatserna .
därför kommer jag nu att lämna tre kritiska synpunkter som tycks oss behöva höras om vi verkligen vill , inte bara i ord utan i sak , &quot; utforma det nya europa &quot; för att använda den ambitiösa titeln på kommissionens dokument och prodis tal .
den första kritiska synpunkten , och i mina ögon den allvarligaste , åsyftar en viss tendens till en litet storvulen självförnöjelse från kommissionens sida när det gäller europeiska unionen själv och en summarisk och rent av nedlåtande syn på våra partner .
en perfekt demonstration på denna frånstötande last finns i de första raderna i kommissionens meddelande .
man talar där om europeiska unionen såsom &quot; ett levande bevis på att fred , stabilitet , frihet och välfärd kan ges åt en världsdel och såsom en modell för hela världen som visar den rätta vägen framåt &quot; innan den avslutar med &quot; att våra grannar har möjlighet att ansluta sig till denna välfärd och att vi har ett drömtillfälle för att göra det möjligt för dem &quot; .
jag tror att en mer nyanserad och sträng diagnostik skulle vara på sin plats .
den idé enligt vilken euron skulle ha främjat ett samförstånd om återhållsamma löner verkar dessutom inte bekräftas av europeiska centralbankens nervösa och upprepade ålägganden till facken , som bedöms vara alltför krävande .
min andra kritik utgår egentligen från den första .
denna extrema svårighet att se verkligheten i sina motsägelser och , i detta fall , att än en gång ifrågasätta sig själv ligger bakom de allvarliga begränsningar som så lägligt anges av prodi , av viljan att bemöta medborgarnas krav .
till exempel åtminstone vad gäller de länder som jag känner väl , tvivlar jag på att den avsikt , som upprepas tre eller fyra gånger i kommissionens dokument , att , jag citerar , &quot; reformera systemen för social trygghet , hälsovård och pension i europa i ett sammanhang av inbesparingar av offentliga utgifter &quot; bemöter de personers förväntningar vars förtroende vi säger att vi vill återvinna .
min tredje kritik är resultatet av de båda iakttagelserna : den svaga diagnosen och låsningarna på vägen till de nödvändiga förändringarna leder till ett projekt som verkar omfattas av ett svårt handikapp på grund av mångfalden av allmänna idéer , en litet impulsiv metod och därmed också av brist på uthållighet .
men ingenting är förlorat .
det handlar om en utgångspunkt , vi har fem år på oss för att lyckas , i den mån den politiska viljan finns och uttrycks med tillräcklig kraft och tydlighet .
min grupp är för sin del fullt ut besluten att bidra till det .
fru talman ! att reformera och demokratisera europeiska unionens institutioner är avgörande för den historiska och moraliska utmaningen om utvidgningsprocessen .
detta var öppningsanförandet av kommissionens ordförande , prodi , när han presenterade europeiska kommissionens strategiska mål för de kommande fem åren .
vi väntar på vitboken om europeiska unionens förvaltning och avvägningen mellan medlemsstaternas regeringar och europeiska unionens institutioner som skall offentliggöras i sommar .
i denna speciella fråga anser jag det viktigt att vi tar upp reformen av kommissionens interna beslutsprocesser .
kommissionen har i sitt förslag till den förestående regeringskonferensen angivit att den föredrar att se mindre medlemsstater förlora sin automatiska rätt att nominera en ledamot till europeiska kommissionen .
detta gäller ett scenario där europeiska unionen har över 25 medlemsstater som medlemmar .
jag vill verkligen inte se en europeisk union byggas i två skikt .
jag anser att detta skulle strida mot romfördragets anda och syfte och alla andra senare fördrag .
det måste finnas likställdhet vad gäller nationell representation inom kommissionen och inom alla andra europeiska institutioner .
jag vill påminna dem som strävar efter att ta bort rätten för små medlemsstater att nominera en europeisk kommissionär att usa ger små stater samma erkännande som större stater i förenta staternas senat .
nästan var och en av de 50 staterna i usa har två valda ledamöter i förenta staternas senat , oavsett dess befolkningssiffra .
varje framtida reform av europeiska unionens fördrag kommer at kräva en folkomröstning i mitt land .
det skulle bli mycket svårt för dem som föreslår en &quot; ja &quot; röst för ett sådant framtida fördrag att få stöd av det irländska folket , om vi förlorar vår rätt till vår kandidat till europeiska kommissionen .
otvivelaktigt skall reformeringen av europeiska rådet också innefattas i denna vitbok om europeiska unionens förvaltning som skall offentliggöras i sommar .
återigen finns speciella politikområden som borde falla under de nationella medlemsstaternas ansvar .
jag tror inte att det finns ett brett stöd i europa för att införa kvalificerad majoritetsröstning om beskattning , rättskipning och inrikes- och utrikesfrågor på europeiska unionens nivå .
enligt artikel 99 i romfördraget måste beslut fattade på eu-nivå om skatteändringar för närvarande vara enhälliga .
jag anser att detta förslag bör kvarstå då en generell europeisk beskattningskod skulle försämra snarare än öka europeiska unionens verksamhet .
jag stöder utvidgningen av europeiska unionen .
jag stöder institutionella förändringar för att kunna garantera att utvidgningen av unionen sker på ett effektivt och strukturerat sätt .
vi måste emellertid komma ihåg att den allmänna opinionen på 370 miljoner människor i den europeiska unionen är en viktig faktor då man förändrar eu-fördragen .
förändringar bör inte ske alltför snabbt och får inte vara alltför vittgående , i annat fall kommer den allmänna opinionen att göra en ratificering av varje framtida eu-fördrag mycket svår att få igenom .
fru talman ! jag skall tala för de radikala italienska ledamöterna .
herr ordförande i kommissionen , ni sade nyss att inga politiska instanser upprättar femårsplaner .
detta är sant om vi tänker på rysslands planer på trettiotalet , men ni meddelade själv för några månader sedan , när er mandatperiod började , för talmanskonferensen att ni faktiskt skulle lägga fram ett program för mandatperioden , det vill säga de stora linjerna för den europeiska regering ni leder och vars verksamhet vi ägnar oss åt i dag .
om det nu än skall vara ett regeringsprogram eller ett tendentiöst program ger en analys av det dokument ni har överlämnat till oss och det tal som åtföljde det inte annat än en katalog över goda avsikter eller snarare över frågor som är på tapeten , utan att man får intrycket att kommissionen tar klar ställning i någon av dessa frågor , det vill säga utför den uppgift som tillkommer europeiska kommissionen .
i detta parlaments kammare har vi tidigare upplevt stora debatter om stora strategiska val som kommissionen har framfört , i kraft av sin initiativrätt , mer som ballon d &apos; essai , som förslag som sedan har rönt mer eller mindre framgång , men som ändå har bidragit till att europeiska unionen har integrerats och utvecklats .
i detta fall har vi verkligen ett antal budord , herr ordförande : man räknar upp en hel rad frågor men ger , om ni tillåter , intrycket att kommissionen inte på någon punkt på något sätt vågar säga &quot; i fråga om detta skulle vi behöva göra så här &quot; .
jag tycker bara ni verkligen tryckte - för mycket tycker jag - på en punkt , det vill säga på att den uppgift ni ser som den nästan högst prioriterade är att avveckla &quot; onödig &quot; verksamhet .
låt oss emellertid se upp , herr ordförande , för vi har haft en förtroendekris för kommissionen och vi har satsat på den här kommissionen - åtminstone har en majoritet av detta parlament satsat på den här kommissionen - just för att reformeringen av kommissionen framför allt skulle innebära en förstärkning , en ny identitet , en ny medvetenhet om att åter ledas av en säker hand .
låt oss tänka oss att kommissionen skulle vilja avveckla eller skulle erbjuda sig att avveckla till exempel de befogenheter den har fått genom fördragen , att verkställa den gemensamma politiken , eftersom den inte tyckte sig vara kapabel till detta .
vad är det vi begär av en regering ?
vad begär vi av denna tvetydiga och speciella så kallade struktur , europeiska gemenskaperna ?
det är bra att de gemensamma resurserna har en övernationell regering och att de inte delegeras till medlemsstaterna eller kontoren för tekniskt bistånd ( bat ) , vilket har hänt tidigare .
ni verkar föreslå oss samma meny men på ett sämre sätt , eftersom ni som ni säger begränsar er till uppgiften att skapa någon vitbok , som ni erbjöd oss .
det jag fruktar - även om ni skakar på huvudet , herr ordförande - är att detta betyder det som vissa länder tycker sedan många år , det vill säga att kommissionen skall vara ett bra sekretariat till ministerrådet .
om det är denna roll kommissionen avser att spela under de kommande fem åren är vi , som är övertygade federalister , säkra på att detta inte är rätt väg att gå och vad detta beträffar kommer vi att ställa er till svars och bedöma vad kommissionen har för avsikt att göra .
reformen är viktig men om den leder till en kantstött kommission , till att dess övernationella befogenheter reduceras och försvagas , handlar det om systemet för den europeiska integrationen , det som grundarna skapade för europeiska kommissionen .
vad de andra punkterna beträffar , herr ordförande , tar jag den om ekonomisk politik och socialpolitik som exempel : visst befinner sig den europeiska sociala modellen i djup kris , visst är arbetslöshetsproblemet det främsta problemet som inga av våra politiska åtgärder har lyckats lösa - och inte av en tillfällighet , men det är inte så att det kan lösas genom att man sammanställer den problemlista vi talade om tidigare , utan att ha en klar vision , ett förslag , det som gör att det finns ekonomier i vårt europa vars takter hör till de snabbaste och som - inte av en tillfällighet - är de ekonomier som har förstått att sätta en flexibel arbetsmarknad och industri som främsta mål .
om vi fortsätter att trassla in oss i förslag som hittills har burit mycket dålig frukt vet jag inte hur vi skulle kunna göra och vad kommissionen kan göra .
detsamma gäller utvidgningen som självändamål , utan att den hänger samman med en mycket mer effektiv reform av europeiska unionen och dess strukturer , med förslag som kommissionen lika gärna skulle ha kunnat framföra vid regeringskonferensen .
herr ordförande , jag vill säga er någonting positivt , kanske tvärtemot somliga kollegers åsikt , vad beträffar det telegram ni skickade till den österrikiska regeringen .
ert ställningstagande övertygade oss : ni gjorde rätt i att inte ytterligare isolera detta land .
fast sedan får vi i handling se vilka de konkreta gesterna blir .
herr ordförande , jag upprepar : det är en vision som enligt vår mening är något närsynt .
framför allt saknas initiativ på de områden jag har tagit upp , till exempel vad gäller balkan .
är det möjligt att fortsätta att hålla balkan utanför utvidgningen , utan att tycka att kroatien , makedonien och andra länder även de har rätt att vistas i detta gemensamma hus ?
fru talman , herr prodi ! jag vill gärna berömma ert förslag om en genomgripande decentralisering av unionens verksamhet och fråga varför ni i så fall lägger fram en förteckning över lagar som är centraliserande .
jag minns er företrädares tal för fem år sedan .
han lovade precis som ni &quot; mindre och bättre &quot; , men santer slutade med att ha levererat &quot; mycket mer och mycket sämre &quot; , och jag tror inte att ni heller kan leverera den utlovade varan .
ni talar om en decentralisering , men centraliserar .
förteckningen över lagar är ju en lång uppräkning av frågor där medborgarna förlorar inflytande och där ni , herr prodi , tar bort detta från medborgarna t.o.m. när det gäller sociala frågor .
ni talar om större öppenhet , men lägger fram förslag som sekretessbelägger handlingar som i dag inte är det .
er kommission är de enda 20 personerna i eu som kan föreslå en minskad lagstiftningsmängd .
det kan inga lokala politiker när man först har lagstiftat i bryssel .
lagkatalogen från kommissionen bör därför åtminstone åtföljas av en lika stor katalog över uppgifter som återsänds till medlemsstaterna och medborgarnas demokrati .
annars växer ju lagmängden ständigt i bryssel .
vi har passerat 10 000 lagar och lika många lagändringar och ansökarländerna har fått 26 000 handlingar skickade till sig , som i det polska parlamentets behandling motsvarar 140 000 sidor .
det är alldeles , alldeles , alldeles för mycket redan i dag .
bryssel skall bestämma mindre och överlämna fler beslut till medborgarna , regionerna och medlemsstaterna , och de beslut som blir över skall endast handla om gränsöverskridande frågor som de nationella parlamenten inte längre kan besluta om på ett effektivt sätt .
och arbetet i bryssel skall ha en mycket högre kvalitet och ske under fullständig öppenhet , så att medborgarna åtminstone kan få litet &quot; medkänsla &quot; när prodi och hans företrädare nu har tagit bort deras rätt till självbestämmande .
till sist bara en kommentar till dell &apos; alba om vad grundarna drömde om : läs de minnen som jean monnet nedtecknat .
det han drömde om var ett litet , praktiskt sekretariat .
det är inte det som prodi är ordförande för i dag .
fru talman ! i morse lade kommissionens ordförande , prodi , fram ambitiösa mål för europeiska unionen för de kommande fem åren , verkligen lovvärda mål , för att skapa en stark och effektiv europeisk närvaro kännbar i världen : framgång med utvidgning , klara utmaningen att sälja e-europa och införa bättre förvaltningsprinciper .
vi godtar att européer , i synnerhet den yngre generationen , måste ges ett brett perspektiv på var europa kommer att befinna sig under kommande år .
men hur skall vi lyckas när de tillgängliga resurserna är begränsade och våra institutioners trovärdighet inte är särskilt hög ?
vi måste anpassa denna vision till verkligheten .
här finns tre beståndsdelar som jag skulle vilja lämna som bidrag .
för det första behöver vi en framgångsrik europeisk ekonomi .
vi måste se till att arbetslösheten fortsätter att minska i hela europa , stärka trenden med privatisering och avreglering , uppmuntra till införande av informationsteknik och kunskap om internet , visa att ett elektroniskt europa är ett bra initiativ .
men vi måste undvika att smyga tillbaka till gammalmodig reglering och kväva enskilda initiativ och företagsskapande .
vi får inte vara rädda för globalisering , men vi måste också se till att vi förstår dess politiska effekt på nätverkssamhället .
utan en framgångsrik europeisk ekonomi kan vi inte klara de kommande utmaningarna , framför allt inte utvidgningen .
för det andra måste vi se till att vi lagstiftar enbart när så krävs - subsidiaritet .
göra mindre men bättre - en central politisk punkt hos den senaste kommissionen - måste vara målsättningen även för denna kommission .
vi kommer att granska detta noggrant när vi skall utforma de årliga programmen om förslag till lagstiftning .
bonde hade rätt när han sade att det finns denna föreställning om att göra mindre men bättre , och sedan får vi plötsligt se ett årligt program för år 2000 med 500 förslag och rekommendationer som verkar gå mot olika mål .
vi måste bestämma vad som skall prioriteras och säkerställa att man får valuta för pengarna i vart och ett av dessa program .
till sist måste vi se till att det blir en verklig och genuin reform av europeiska kommissionen .
ja , kommissionen - fördragens väktare - är avsedd att vara ett oberoende organ men det måste även vara ansvarigt inför europeiska medborgare genom vårt parlament .
det informationsproblem som bonde just nämnde behandlas som ett tecken på att kommissionen verkar begränsa informationen till oss , som medborgare och som parlamentariker , fastän vi har rätt till den enligt fördragen .
kommissionen är egentligen inte i dag en europeisk regering .
kommissionen avspeglar inte majoriteten i detta speciella parlament .
vi i parlamentet har en stor roll att spela för att utforma förvaltningen i europa .
denna elektroniska förvaltning måste därför vara en lyhörd förvaltning så att vi faktiskt kan arbeta tillsammans och inse att var och en av institutionerna i europeiska unionen har sin tillämpliga roll att spela .
därför behöver vi trovärdighet , sammanhållning och tillförsikt om att vi genom att arbeta tillsammans kan återställa våra medborgares bild av europeiska unionen .
fru talman , herr kommissionsordförande ! jag samtycker fullt ut med tankarna i de förslag som gjorts av min kollega heidi hautala vad gäller kommissionens strategiska mål för de kommande fem åren .
jag kommer för min del att hålla mig till ett ämne som ni inte har tagit upp och som hade planerats och gäller kommissionens arbetsprogram för år 2000 .
jag är medveten om budgetårets begränsningar eftersom vi arbetar inom ramen för det aktuella fördraget och är begränsade av dess funktionsregler - jag tänker särskilt på en viktig fråga som är skattefrågor .
men jag skulle faktiskt inte vilja tala om skattefrågor .
jag kommer att börja med att välkomna vissa förslag som ni lägger fram inför programmet för år 2000 .
jag tänker på alla förslag i fråga om livsmedelssäkerhet som är ambitiösa och viktiga och jag tänker också på sjösäkerhet efter de båda oljeutsläppen utanför bretagnes kust och i turkiet .
det är bra att kommissionen reagerar snabbt i det avseendet .
när det gäller andra frågor anser jag däremot att man skulle kunna vara mer ambitiös och gå snabbare .
och jag skulle vilja lämna ett antal positiva förslag , där tänker jag framför allt på det sociala området , miljön och uppföljningen av seattle .
en inledande anmärkning : ni sade att det är nödvändigt att åter försona de europeiska medborgarna med deras institutioner , något som är självklart , och jag tror således att det är viktigt att vi undrar över vad som i främsta ledet upptar medborgarnas tankar .
jag tror till exempel att på det sociala området räcker det inte med att utfärda ett meddelande om ett program för sociala åtgärder .
det måste gå snabbare .
ni måste lägga fram ett nytt program för sociala åtgärder för oss i slutet av året .
en fråga , slutligen , som har ingått i de senaste nyheterna och fortfarande upptar en stor plats i dem är frågan om företagsnedläggning och kollektiva uppsägningar .
vi arbetar på grundval av ett aktuellt direktiv som har visat sig ha sina begränsningar och vi skulle vilja - och jag ger er ett förslag - se över denna direktivtext så att vi får ett effektivare direktiv vad gäller sysselsättningsskydd och också effektivare vad gäller eventuella sanktioner mot dem som inte följer texten .
när det gäller miljön aviserar ni ett förslag till beslut om ett sjätte åtgärdsprogram om miljö och det är mycket bra .
man har sagt mig - men ni skall kanske dementera mina uttalanden - att det inte finns några exakta mål och någon tidsplan för genomförande i den text som ni skall föreslå oss .
jag tror personligen att det är nödvändigt att ha beräknade mål och en verklig tidsplan för genomförande .
jag tror också att när det gäller frågan om enskilt ansvar är det glädjande att vi äntligen har en vitbok , jag talar då om enskilt ansvar gentemot miljön , men jag vill påminna om att parlamentet har begärt ett lagstiftningsinitiativ i sex år , och att vitboken naturligtvis aviserar en sådan lagstiftning , men när ?
där vill jag också uppmärksamma er på att processen måste påskyndas .
slutligen den sista delen , efter kyoto skulle det ändå vara sunt om vi skulle snabbt komma fram till exakta förslag och jag vill sluta med att säga ett ord om wto .
jag tror att tanken på att åter sätta i gång en ny global period inte är en dålig tanke men jag tror och upprepar att först måste verkligen kommissionen ge oss förslag för att ändra wto : s funktionsregler .
kommissionen har en inre roll , men också en roll i världen .
det verkar som om europeiska unionen bör ligga till grund för en omvärdering av wto : s funktionssätt , en omvärdering som bör leda till att vi ger exakta förslag i stadgehänseende .
fru talman ! ni talade om grundläggande politiska värderingar och en av de grundläggande politiska värderingarna , till och med mer grundläggande än demokratin , är respekten för andra .
därför anser vi att ni gjorde rätt i att skicka ett meddelande , och att de som kritiserar det kanske fortfarande lider av sviterna av en bolsjevitisk eller nazistisk kultur , för demokrati innebär att föra en dialog med andra och låta dem förstå när de felar , men också lyssna på deras skäl .
att utvidga får inte innebära att urvattna , det vill säga det får inte innebära att man utvidgar riskerna . detta har nationella alliansen upprepat i tio år i denna kammare .
kandidatländernas förhoppningar är minst lika viktiga som våra nuvarande medborgares förhoppningar , vilka börjar bli allvarligt besvikna på hur detta europa fungerar när man inte löser de viktigaste problemen .
utvidgningen kräver alltså stränghet , att man respekterar de villkor som - om det blir nödvändigt - bör omformuleras vad vissa grundläggande frågor beträffar : det som har hänt i rumänien , med konsekvenser ända till belgrad - den ekologiska tragedin - men framför allt att likgiltigheten inför de stora säkerhetsproblemen fortsätter att breda ut sig .
än i dag finns inga slutgiltiga lösningar för kontroll över kärnkraftverken i östrepublikerna .
man måste alltså ha resurser att spendera innan man går vidare mot en utvidgning , för att äntligen skapa en europeisk kontrollstyrka med uppgift att övervaka kvalitet och driftsförhållanden för att skapa en ny värld där vissa tragedier inte längre hör hemma .
jag skulle också vilja säga några ord om afrika , fru talman .
den tredje och fjärde världen är övergivna : det skulle räcka med en dollar , en och en halv euro , för att rädda många barn .
europa som är så demokratiskt , som är så progressivt , tiger och tar inte på sig dessa tragiska problem , under tiden som halva afrika dör i aids och andra sjukdomar .
ett sista påpekande om internet och globaliseringen .
globaliseringen av ekonomin får inte bli en likriktning av produkter och kvaliteter , liksom globaliseringen av politiken inte får bli en utslätning av värderingar , av förhoppningar , av entusiasmen .
de folk som inte deltar , och som sakta drar sig undan , ger utrymme för en oligarki som tar makten och lämnar kontrollen till ett fåtal .
vad internet beträffar : europa måste äntligen ha modet att säga att det krävs regler .
tillåt mig här att , som privatperson , applådera de pirater som genom att handla som de gör tvingar världen att fundera över det enda system som inte har några regler i dag .
vi är en reglernas värld : låt oss ge även internet regler och på så sätt ge medborgarnas framtid regler och hopp .
fru talman ! som skattebetalare i padanien har jag redan känt av uttaxeraren prodis bett på den tiden då han var regeringschef i italien som padanien också skattemässigt är underställt .
jag blev bekymrad när jag lyssnade på honom nu när han antydde nya resurser , ett koncept som lätt kan översättas med nya skatter och pålagor bland annat inför utvidgningen , det vill säga att nya stater träder in i unionen .
men varför betalar inte de sin inträdesbiljett själva ?
mina padanska väljare som tack vare prodi redan har betalat det som i italien går under namnet europaskatt - som bara delvis har återbetalats - har absolut inte för avsikt att , fortfarande tack vare prodi , betala en skatt till för någon annan .
fru talman , herr kommissionsordförande , ledamöter av kommissionen ! fem månader efter sitt tillträde har kommissionen angivit i vilken riktning den vill styra europeiska unionen .
det har blivit en ambitiös men även högtravande handling .
är det inte patetiskt att säga att &quot; världen ser upp till europa &quot; ?
dessutom är världsdelen europa så mycket mer än de femton medlemsstaterna i europeiska unionen .
garanterandet av fred , demokrati och mänskliga rättigheter i , märk väl , hela europa är att sikta litet väl högt .
jag är väldigt nyfiken på hur kommissionen tänker förverkliga det här .
den europeiska integrationsmodellen som en rik källa för världsstyre , är det detsamma som export av storskalighet och maktkoncentration ?
kommissionen anser att utrikespolitiken kan lyckas om var och en vet exakt vem som styr !
vem är det då ?
hela kommissionen , dess ordförande kanske , rådet ?
för den nya ledningen av europa behövs starka institutioner , säger ni , medan kommissionen samtidigt vill koncentrera sig på sina kärnuppgifter .
det senare håller vi gärna med om .
det är verkligen hög tid att institutionerna inskränker sig till problem som verkligen är gränsöverskridande och slutar smycka den europeiska vagnen med befogenheter som tagits från de nationella myndigheterna .
vid flera tillfällen i texten talas det om gemensamma värden .
tyvärr saknar jag en hänvisning till de normer som hör dit .
man kan undra var de normerna och värdena är hämtade från .
jag är övertygad om att bibeln , guds ord , är den enda rena källan till goda normer och äkta värden .
den insikten är en viktig del av traditionen i vår världsdel och den förtjänar att bli erkänd
fru talman , herr kommissionsordförande , mina damer och herrar ! jag vet inte vad jag skall hålla mig till - de strategiska målen för perioden 2000-2005 eller till ert tal om perioden 2000-2010 ?
har ni redan inkluderat er andra mandatperiod ?
men , allvarligt talat .
unionen som håller på att utvidgas behöver stärkas genom bantning och begränsning .
för det första , bantningen .
det ni säger i ert program om att koncentrera sig på kommissionens kärnfrågor är bara en första början .
hela unionens verksamhet måste föras tillbaka till politikens kärnområden .
de omfattar marknadens sociala och ekologiska inriktning , säkrandet av valutan , garantin för de medborgerliga rättigheterna inom unionen och företrädandet av de gemensamma intressena utåt .
här gäller det inte bara att tala med en röst i världen , utan det handlar snarare om vad vi vill säga med denna röst .
för det andra heter det nya modeordet flexibilitet .
men en tilltagande flexibilisering kan bli eller hotar mycket snabbt att bli till ett samarbete på regeringsnivå .
vi måste benhårt hålla fast vid sammanhållningen av medlemsstaterna med hjälp av gemensamma beslutsorgan .
det gäller för övrigt också för införlivandet av det civila samhället , som kan betraktas som positiv .
men medborgarna behöver inga nya organ eller institutioner och absolut inte någon ny sammanblandning av ansvarsområden .
öppenhet betyder inte större tillgång till mer papper , utan öppenhet för medborgarna är att äntligen få mer klarhet om vem som beslutar när och med vilket berättigande i bryssel och strasbourg .
det är öppenhet !
för det tredje kan och får europeiska unionen inte utvidgas gränslöst .
dess gränser bestäms inte av hur många stater som vill vara med , utan av hur många stater som den klarar av .
om priset för utvidgningen vore en uppmjukning eller rent av en upplösning av den befintliga unionen , då får man inte betala det priset .
det skulle vara för högt , för övrigt inte bara för dess medlemsstater , utan också för de stater som vill bli medlemmar i unionen .
en union enbart som ett geostrategiskt koncept har inte någon framtid , lika litet som en union som enbart är en frihandelszon .
men unionen förblir något mer än en marknad och får sin legitimitet av europas folk enbart om den uppfattar sig som en ödesgemenskap .
detta är långt mer än enbart er nya ekonomiska och socialpolitiska agenda eller en ny och bättre livskvalitet .
inte bara kommissionen , inte bara europaparlamentet , utan också folken och staterna i vår europeiska union måste finna nya svar på frågan hur och för vad vi vill leva och agera gemensamt .
här handlar det inte om något mindre än att uppfinna europeiska unionen på nytt , utan att förstöra det som redan existerar !
herr talman ! enligt europeiska liberala och demokratiska partiets grupp är kommissionens och hela unionens viktigaste uppgift under de närmaste åren att genomföra utvidgningen med framgång .
kommissionen skall i förhandlingarna målmedvetet sträva efter att varje ansökarland skall kunna gå med i unionen snarast möjligt .
å andra sidan måste man se till att inte omintetgöra hittills uppnådda resultat eller målsättningarna för integrationen .
för att undvika detta har den liberala gruppen framfört ett önskemål om att man vid regeringskonferensen skall överväga olika modeller för en differentierad integrering och att man skapar en koncentrisk union med en federationskärna och en mindre integrerad yttre cirkel .
det är uppenbart att unionens interna differentiering tas upp på regeringskonferensen .
behandlingen av denna fråga kräver fördomsfrihet .
det räcker inte med att tekniskt förbättra det flexibla samarbetet , utan man måste också diskutera utvecklingen av de egna institutionerna för avant garde-länderna , såsom bland annat jacques delors har föreslagit .
på detta sätt kan vi skapa en ännu effektivare , tydligare och mera demokratisk beslutsprocess .
jag hoppas att komissionen lämnar ett eget förslag till hur den institutionella och övriga differentieringen i den utvidgande unionen bör genomföras .
fru talman , herr kommissionsordförande , mina damer och herrar ! ert inspirerande anförande , herr prodi , har förfört mig .
det väcker förväntningar men det kan också leda till besvikelse .
det har att göra med det som van velzen sade alldeles nyss , med skillnaden mellan ord och handling .
unionens utvidgning kommer sig av vår längtan efter fred , säkerhet och stabilitet .
ni vill lugna de nya staterna och även den europeiska opinionen .
vi ser dock med våra egna ögon att det motsatta sker i dag .
vi ser hur rädslan och oron ökar , även i de områden där arbetslösheten inte är hög och välfärden är väldigt stor .
vi måste kunna ge våra medborgare en hemkänsla , sade swoboda , och det har han rätt i .
det är en plats där vi alla delar samma värden och där var och en har sin uppgift och sitt ansvar .
det har antagligen att göra med de normer som van dam talade om .
det är nämligen subsidiaritet . tydligt ansvar för alla ledningsnivåer , partner och inte konkurrenter i styret .
makten så nära medborgarna som möjligt , där den kan utövas öppet och under insyn och kontrolleras av medborgarna själva .
för det krävs en ny politisk kultur , inte bara i teorin utan även i praktiken , där man tar hänsyn till den verklighet som råder i medlemsstaterna och i regionerna .
regioner som i kulturellt och ekonomiskt avseende ibland är lika viktiga som vissa medlemsstaters intressen .
det nya europa får inte bara utvecklas på bredden utan även på djupet , genom att omsätta våra värden i praktiken och genom ett demokratiskt byggande av en äkta gemenskap .
på det skall kommissionen bedömas .
fru talman , kommissionen lägger idag fram sina strategiska målsättningar för perioden 2000-2005 i form av ett extremt allmänt hållet dokument i vilket de sträva anmärkningarna strukits för att inte alltför mycket såra en del personer .
i den första delen således rörande de nya formerna av europeiskt regerande läser man inte någonstans naturligtvis orden federalism eller superstat .
men det är ändå de som framträder när det är fråga om en stark europeisk institution i vilken enbart de löpande genomförandeverksamheterna decentraliseras och skjuter in sin kollektiva syn i en oklar enhet där regeringar och nationella parlament är beblandade med regionala , och till och med lokala , myndigheter samt med det civila samhället , samtliga utsedda , utan någon hierarkisering såsom , jag citerar : &quot; deltagande part i europeiska frågor &quot; .
dessa tvetydigheter döljer många missuppfattningar och främst om våra värderingar .
det räcker nämligen inte med att åberopa demokrati för att vara demokrat .
man måste framför allt acceptera att medborgarna fritt fattar beslut på den nivå där de objektiva villkoren för en nära , lojal och öppen demokratisk debatt bäst finns samlade , det vill säga huvudsakligen på nationell nivå .
kommissionens meddelande i sin helhet är emellertid just uppbyggt på motsatt påstående enligt vilket det skulle vara nödvändigt att under förevändning att bättre försvara folket fortsätta att begränsa deras marginal för självständigt val ytterligare genom nya föreskrifter , nytt införlivande av politik eller nya tvingande rättsliga strukturer såsom förslaget till stadga om så , felaktigt , kallade grundläggande rättigheter .
jag betonar &quot; felaktigt &quot; eftersom den i själva verket skall minska dessa rättigheter .
i gruppen unionen för nationernas europa är principerna mycket annorlunda .
vi vill försvara europas länder men också respektera folkens val .
det är inte alls cirkelns fyrkant .
vi måste nämligen överge de omoderna federalistiska modellerna , de modeller som satts upp av dem vars idéer om europafrågan härrör från jean monnets memoarer .
vi måste tvärtom öppna de europeiska institutionerna för den moderna världen genom att uppfinna en dynamik av variabel geometri som respekterar nationerna .
detta är den stora idén om ett nytt ledningssätt som vi skulle ha velat finna i ert meddelande , herr ordförande . tyvärr fanns det inte där .
fru talman , herr kommissionsordförande ! ni påstår att ni utformar ett nytt europa men ni saknar tyvärr en väsentlig förutsättning : förtroende .
man kan nämligen inte dra till sig miljoner européers förtroende när man inte är värd det .
och hur skulle ni kunna vara värd ett förtroende efter galna ko-affären och santer-kommissionens avgång på grund av korruption ?
ni bär ansvaret för miljoner arbetslösa och miljoner fattiga samt ökande utsatthet och nöd på grund av er extrema handelsutbytespolitik och ultraliberala politik och på grund av tvångsmarschen till den gemensamma valutan .
ni har velat ha och har ordnat avlägsnandet av de inre gränserna och ni har sålunda utsatt europa för en explosion av kriminalitet och osäkerhet och en flodvåg av okontrollerad invandring .
ni föreslår nu att en handfull tjänstemän skall få hela beslutandemakten och göra staterna , de lokala myndigheterna och de icke-statliga organisationerna , där alla för övrigt har lika villkor i sitt beroende till bryssel , till enkla verkställare av beslut som kommer ovanifrån .
i ert fjortonsidiga dokument nämns inte en enda gång de nationella parlamenten , som likväl i motsats till kommissionen består av folkvalda ledamöter .
men de har visserligen inte någon roll i er strategi .
ni vågar inte ens kalla saker och ting med sitt rätta namn och ni gömmer er bakom en låtsad inne-semantik genom att kalla det för &quot; guvenörskap &quot; , det som inte är något annat än en federal enväldig centralregering .
efter att i åratal ha försökt övertyga genom att tala om delad suveränitet medger ni nu ert yttersta mål : att sälja ut den europeiska suveräniteten , vare sig den är nationell eller lokal , till en världsregering i vilken ni inte ens hoppas på att få en avgörande plats .
ni vågar slutligen fördöma och sanktionera , eller låta fördöma och sanktionera , miljoner österrikares fria och demokratiska val av det skälet att ni inte tycker om resultatet .
och på samma gång stöder ni det kommunistiska kina och har handel med länder som öppet bryter mot mänskliga rättigheter sedan årtionden tillbaka .
i dag igen går de europeiska parlamentsledamöterna angrepp mot ett telegram från prodi till kansler schüssel som likväl påtagligen inte är en sympatiyttring utan en politisk manöver .
ert skryt bedrar inte någon eftersom , och det vet ni mycket väl , vare sig ni vill eller inte behöver ni österrike för att reformera fördragen och harmonisera skattesystemet för sparande .
ni använder österrike som en bekväm fågelskrämma .
era kommissionärer är förvisso inte de enda som är ansvariga .
de regeringar som stöder er av slapphet eller av ideologiska skäl är det också .
bryssel är inte vi alla som ni påstår , utan det är ni alla .
ljug inte mer , ni struntar väl i vad europas folk vill .
européerna är bara fria att välja mellan er bästa av världar och att ställas vid skampålen .
mer än tio år efter sovjetunionens upplösning osar era förslag av gulag med tillägg av en lenande moralism .
vi var en del av den lilla klick som pekade ut den kommunistiska diktaturen .
vi är och kommer att förbli bland dem som bekämpar en europeistisk diktatur och vi uppmanar alla europas folk att gå med i motståndet mot era ohyggliga förslag .
de europeiska demokratiernas räddning finns i staten såsom nation och i den nationella staten och europas räddning finns i samarbetet mellan nationerna i europa .
( några applåder )
ordförande prodi , ni har i dag presenterat ett femårsprogram för kommissionen med många mål som man kan instämma i , ett program som består av scenarier och ledmotiv , och det är därför riktigt att hålla sig kvar vid de stora dragen , bortom de konkreta inslagen .
av era ord och det dokument ni har överlämnat till oss verkar det som om en fråga som ligger er , herr ordförande , och mig varmt om hjärtat har hamnat i skymundan : solidariteten , inte så mycket på det internationella planet som internt .
ärkebiskopen i milano , hans högvärdighet carlo maria martini , uppmanar alla politiker och särskilt sådana som ni och jag , herr ordförande , sådana som kulturellt och värdemässigt grundar sitt politiska engagemang på katolicismen , att omvärdera en utvecklingsfråga som förutom den ekonomiska vinsten mycket , oerhört mycket , berör dem som har det sämst ställt , de utstötta .
det är en stor fråga , den om de som har det sämst ställt , en stor fråga som påminner oss om hur svårt och komplicerat det är att fastställa mått på framsteg och hur otillräckligt det är att bara se till inkomsten per capita .
det påminner oss också om behovet av en ny utvecklingsmodell som är stadigt förankrad i en kultur med socialt engagerade katoliker , vilka betraktar det civila samhället , de samhälleliga instanser som allmänheten främjar och understöder , som de sundaste instrumenten för att bygga solidaritet .
på så sätt betonas den grundläggande elementet för varje individs utveckling : hennes frihet , som kommer före den ekonomiska vinsten .
denna samhälleliga frihet som yttrar sig i initiativ till förmån för dem som har det sämst ställt ger återbetalning i form av rättvisa och samhällelig balans .
herr ordförande , de offentliga institutionerna skall inte bara följa ekonomiska kriterier .
de måste rikta in sig på service till individerna och arbetet med att bygga upp var och ens frihet , naturligtvis utan att glömma att allt detta inte får och inte skall stå i motsats till behovet av att skapa företagsamhet , att investera och riskera . i ett ordentligt och målinriktat system kan entreprenörerna bidra till samhällets tillväxt och till solidariteten i betydande omfattning .
i globaliseringens tidevarv , globaliseringen som vi dock vill ge en ram av fasta regler som ger de ekonomiska aktörerna och konsumenterna trygghet , får inte europeiska kommissionen glömma solidariteten och betona att den skall tillämpas i alla medmänskliga relationer .
vår historia har lärt oss att hjärtat måste finnas med i politiken .
vi hoppas att vitboken och era och kommissionens handlingar kommer att visa detta i praktiken .
fru talman , kommissionsordförande , kolleger ! shaping the new europe är en ambitiös målsättning för kommissionen och för oss alla .
vår ambition och vårt arbete kommer att följas av medborgarna i våra länder , men också av många utanför europa och utanför vår union .
vilken bild får då en intresserad allmänhet och resten av världen av detta femårsprogram ?
mitt svar är : en nystart , en tydligt reformistisk agenda , som bekräftar att 2000-talets union inte vill stanna vid att vara en ekonomisk gemenskap , utan vill vara en värdig gemenskap , som vi tar på allvar .
med rätta säger kommissionen att unionens avsikt är att utveckla och värna om ett solidariskt välfärdssamhälle i globaliseringens tidevarv , ett rättfärdigt och effektivare europa , som också ser sitt ansvar utanför den egna kontinenten utifrån solidaritet och upplyst egenintresse .
vi ser nämligen fattigdom och utanförskap som fredens och frihetens främsta fiende .
med instämmande i vad mina partivänner har sagt och med gillande av grundtonen i ert dokument vill jag rikta uppmärksamheten på två brister , som måste korrigeras i det kommande arbetet .
det första gäller kvinnor , gender eller kvinnors rättigheter .
ni talade om kvinnors medverkan för att öka produktion och tillväxt .
detta är viktigt , men jämställdhet är inte bara nödvändigt för produktiviteten utan också för demokratin i våra samhällen .
det är därför uppseendeväckande att ordet jämställdhet , gender eller kvinna överhuvudtaget inte förekommer någonstans i shaping the new europe .
ni talade om kvinnan i ert tal , men hon nämns inte bland de strategiska målen .
beror detta , herr kommissionär , på att mainstreaming redan är så genomförd i kommissionen att kvinnor inte behöver nämnas ?
hur förklarar ni annars denna frånvaro av kvinnor .
eu får inte bli en union med manligt ansikte .
min andra fråga gäller afrika . inte heller afrika nämns i shaping the new europe , men alla andra kontinenter .
i afrika har vi världens högsta antal flyktingar , världens största samlade fattigdom och en förtärande aidsepidemi .
jag vet att kommissionär nielson och andra gör ett bra jobb , men det krävs att hela kommissionen , också i sina strategiska målsättningar , fokuserar mer på denna kontinent .
slutligen vill jag välkomna kommissionens uttalande och att det i detta för första gången sägs att eu är berett att unilateralt vidta åtgärder till förmån för ökat tillträde till våra marknader för utvecklingsländerna .
min fråga är : när kommer detta att sjösättas ?
fru talman , herr ordförande i kommissionen , ärade ledamöter ! vi har framför oss ett dokument som har avgörande betydelse för europas framtid och öde .
av alla frågorna framträder emellertid direkt två som är intimt förknippade med varandra : freden och stabiliteten i och utanför europa .
det handlar om mål som skall prioriteras .
sedan länge delar vi alla detta synsätt , men vi måste också tydligt hävda att dessa mål inte kan uppnås utan utvidgningen , även om denna skulle medföra kostnader .
i dag är det vår uppgift att för de kommande decennierna välja mellan ett europa som kanske är mindre rikt , men som är en ledstjärna för fred och civilisation för hela vår planet och ett europa som kanske är mer välmående men saknar visioner .
dessa mål kan dock endast uppnås om regeringskonferensen , som kommer att avslutas innan årets slut , ger upphov till en konstitutionell reform som ger kommissionen adekvat och reell makt . kommissionen kan inte fortsätta att bara vara den som verkställer rådets beslut och parlamentets medbeslutande utan måste spela rollen som europas verkliga regering .
parlamentet borde vara den förste att stödja denna reform om det verkligen vill vidga sin roll som uttolkare av européernas vilja och skaffa sig den centrala funktion som tillkommer en union som är sant demokratisk och kraftigt integrerad .
för övrigt kan kommissionen bara ges ansvar för de åtaganden den tar på sig i den utsträckning den reella befogenhet den har medger .
om dessa skisserade möjligheter saknas kommer europa att retirera in i en historia utan framtid .
fru talman , herr kommissionsordförande ! vi kan glädjas åt den globala ambitionen i de angivna målsättningarna , som går parallellt med de utmaningar som europa skall tvingas klara av .
jag noterar att ni anser att berlinmurens fall är den väsentliga faktorn i sekelslutet .
denna händelse bör leda till utvidgning .
jag har lust att snarare tala om återförening än att använda ordet &quot; utvidgning &quot; . det tycks mig ha en politiskt mycket starkare betydelse .
ni återupptar tanken att omcentrera era verksamheter runt de viktigaste uppgifterna och det ingår i målsättningarna för er reform .
i grunden handlar det om att tillämpa subsidiaritetsprincipen .
en klar tillämpning av denna princip kan bara stärka de åtgärder som vidtas och ge medborgarna en klar bild av varje behörighetsnivå .
men , herr prodi , att säga det är en sak men att göra det är en annan !
ni måste således kämpa mot alla institutioners tendens att i allmänhet försöka öka sina befogenheter ytterligare .
jag kommer således att döma efter handling .
under tiden instämmer jag i och uppmuntrar denna tydligt uttryckta vilja i ert meddelande .
två saker är emellertid väsentliga : förenkling och tillämpning av gemenskapsrätten .
1998 var det 123 anhängiggöranden i domstolen på grund av icke-tillämpning eller icke-införlivande av gemenskapsrätten och 25 procent av direktiven om miljöfrågor tillämpas inte eller är inte införlivade .
händelserna de senaste dagarna visar hur nödvändigt det är .
gemenskapsrätten får inte vara utan tillämpning för att den är för komplicerad eller för detaljerad .
unionen får inte falla i den fällan och också i det avseendet beklagar jag att ert meddelande inte går in mer på detaljer .
ni är realistisk i fråga om att välfärdsstaten inte längre kan lösa de problem som uppstår och bland annat arbetslösheten .
jag beklagar dock att ett klart alternativ inte lagts fram .
man borde ha betonat att all understödspolitik förkastas och däremot värderas initiativ och ansvar .
ni framhåller inte åldrandet av befolkningen som kommer att få grundläggande verkningar på vårt samhälles struktur inte bara ur ekonomisk synpunkt utan också på folkhälsoplanet .
det handlar egentligen om en tyst revolution och i det avseendet väntade jag mig mera i ert meddelande .
ni betonar slutligen att den europeiska forskningen står i centrum inför vår framtid .
ni anger emellertid inte vilka medel ni vill sätta in .
de etiska principerna finns också i centrum av denna forskning . i ert meddelande nämns ingenting .
herr ordförande , ni vill ge bättre information till medborgarna . börja då med att stärka banden med parlamentet : vi är dessa medborgares företrädare .
fru talman , ärade ledamöter ! man kan inte annat än instämma i de allmänna linjerna i femårsprogrammet och programmet för år 2000 , som ordförande prodi har beskrivit med sådan glöd i dag .
i de båda dokumenten betonas starkt behovet av att fastställa nya former för europeisk governance och att i detta syfte omvärdera kommissionens uppgifter med stringentare prioriteringar i strävan mot full sysselsättning . detta genom att samordna staternas ekonomiska politik och socialpolitik på ett mer effektivt sätt och - vilket jag tillåter mig att understryka - i första hand de länder som ingår i den monetära unionen och som måste sättas i stånd att utgöra det första exemplet på stärkt samarbete .
i detta syfte nöjer jag mig med att betona tre av de viktiga prioriterade frågor som bör vägleda europeiska unionens verksamhet under de närmaste månaderna , förutom beträffande kommissionens uppgifter också vad gäller att formulera handlingsprogram för unionens regeringar .
för det första att främja och delta i framtagandet av gemensamma projekt för att skapa ett integrerat servicenätverk inom transport- och energisektorerna , med stöd av europeiska investeringsbanken .
för det andra att besluta om investeringar som skall genomföras i de enskilda länderna och via gemenskapens projekt inom de prioriterade sektorerna forskning , innovation och uppvärdering av den mänskliga faktorn , som förpliktelser i åtgärdsprogrammen om sysselsättning .
jag anser att dessa parametrar - särskilt de kvalitativa som är resultat av investeringar i livslångt lärande , fortbildning , anpassningsbarhet och omskolning av de äldsta löntagarna - är mycket mer betydelsefulla och krävande eftersom deras effekter är varaktiga på medellång sikt . de är något annat än bara uppställandet av årliga kvantitativa mål , som alltid kan ifrågasättas , om att skapa sysselsättning eller minska arbetslösheten .
om kommissionen bland annat , vilket även understryks i det portugisiska ordförandeskapets program , kunde verka för en ny fas i den sociala dialogen som är inriktad på en överenskommen strategi för social kompetens och kunskapsspridning , kort sagt en strategi för anställbarhet och en definition av reglerna för den , skulle detta göra det möjligt att ta steget till att löntagarna blir informerade och instämmande deltagare i omstrukturerings- och återanställningsprocesserna .
för det tredje tror jag inte att minskningen av antalet aktiva till följd av att befolkningen åldras är ett oundvikligt öde för europeiska unionen .
inte bara för att det finns marginaler för att öka kvinnors sysselsättningsgrad och för immigration utan därför att man bestämt måste vända den utbredda tendensen till förtidspensionering och att man tidigt drar sig tillbaka från arbetsmarknaden genom att verkligen inte inrikta den samordnade reformen av de sociala trygghetssystemen på betydande minskningar av de framtida pensionsförmånerna utan på att aktivt utnyttja den ökade förväntade livslängden för att förlänga den yrkesverksamma tiden .
fru talman , herr kommissionsordförande , mina damer och herrar ! herr prodi , ni har trätt in full av ambitioner och reformvilja .
såväl ni som era ambitioner är välkomna .
de kommer att behövas för den omfattande uppgift vi står inför .
men för att kunna genomföra alla dessa reformer och driva lagstiftningsprogrammet för år 2001 vidare måste vi vara säkra , inte bara på styrkan hos reformatorn , utan även på de övrigas åsikter .
ni säger att ni inte kommer att dra er för att komma till oss och be om ökade resurser till kommissionen , men kommissionen bör vara medveten om att vi har en begränsad budget att röra oss med .
vi förfogar över 1,27 procent av gemenskapens bni .
inte en euro mer eller mindre .
det kommer inte att vara vi som vägrar dessa nya resurser , ni bör då snarare vända er till rådet .
budgetplanerna är millimeteranpassade .
för att kunna finansiera stabilitetsplanen för balkanländerna måste man förhandla om den så viktiga granskningen av utgiftsområde 4 , och tänk på de svårigheter vi hade med att godkänna budgeten för år 2000 .
jag kan påminna er om att vår politiska grupp , ppe-de , inte tycker om att nya politiska initiativ finansieras på bekostnad av de som redan existerar .
parlamentet och de europeiska ledamöterna bör fastslå de politiska prioriteringarna .
tro inte för ett ögonblick att den budgetreform som ni föreslår kommer att dölja begränsningarna av gemenskapens finanssystem .
det är bra att vi alla i ömsesidigt samförstånd gör en insats för att rationalisera budgeten , men då bör ni vara medveten om att de otillräckliga resurserna , frånvaron av finansiellt självstyre och det bristfälliga genomförandet av budgeten fortsätter att vara angelägna frågor som måste få en lösning .
därför undrar vi : har kommissionen den politiska viljan att lösa dessa ?
fru talman , herr kommissionsordförande , kära kommissionärer , kära kolleger ! strategidokumentet har enligt min åsikt två tydliga svagheter .
det hjälper inte att författa en ny ekonomisk och social agenda , när man inte har arbetat av den gamla .
jag talar om transportpolitiken eller om regionalpolitiken .
för båda områdena har ni med kollegerna palacio och barnier utmärkta kommissionärer , och trots detta tillmäter ni dessa områden för liten betydelse i ert strategidokument .
beträffande transportpolitiken är det viktigt att denna utformas ekonomiskt och miljöpolitiskt förnuftigt i europeiska unionen , och detta innan andra stater ansluts .
om kommissionsordföranden lyssnade på mig , så vore jag tacksam , men det är ju inte nödvändigt .
jag ger er tre exempel på detta .
för det första : vi behöver en förnuftig avreglering inom järnvägssektorn , ty vi vill föra över godstransporterna från vägarna till järnvägarna .
det är ekonomiskt och miljöpolitiskt klokt .
utan avreglering kan vi inte åstadkomma någon förnuftig transportpolitik .
samma sak gäller den europeiska flygsäkerheten .
medborgarna har inte någon förståelse för att vi avreglerar lufttransporterna , medan det i luften finns kvar 15 olika sektorer , som kontrolleras nationellt , som medför ekonomiska nackdelar för flyglinjerna och som förstör miljön .
här måste ni också beta av er föredragningslista .
herr kommissionär ! regionalpolitiken nämns alltför litet i ert dokument .
den sociala och ekonomiska sammanhållningen inom eu är en avgörande uppgift för denna gemenskap .
om vi inte åstadkommer den , kommer medborgarna i de missgynnade områdena också att vara rädda för utvidgningen .
vi måste klargöra för dem att vi kommer att använda de närmaste fem åren till att stödja de missgynnade områdena och med en klok användning av medlen göra dem till rika områden .
då är även de beredda att verkligen rösta för en utvidgning och vara med om att genomföra den .
herr kommissionsordförande ! om vi inte lyckas åstadkomma en uttalad solidaritet mellan de rika och fattiga regionerna , då kommer denna union att bli fattigare , och den kommer inte att finna något bifall hos befolkningen !
herr talman , herr kommissionsordförande , värderade kommissionärer , värderade kolleger ! när vi utformar nya program , får vi inte glömma de äldre program som håller på att genomföras .
med tanke på detta är det bra att kommissionens arbetsprogram åter tar upp frågorna i agenda 2000 , den gemensamma jordbrukspolitiken , inklusive fisket , och , för det andra , strukturfondernas verksamhet .
jag hoppas , herr kommissionsordförande , att detta betyder att den pågående omorganisationen av kommissionen inte kommer att skada den mekanism för kontroll och genomförande som finns i agenda 2000 .
frågorna i agenda 2000 gäller naturligtvis ert tredje och fjärde strategiska mål , den ekonomiska och politiska agendan och den högre livskvalitén .
vad man kan utläsa av era texter är i vilken utsträckning de högt ställda målen motsvaras av de resurser som kommissionen avser att ställa till förfogande .
och jag menar inte nödvändigtvis ekonomiska resurser .
för att genomföra agenda 2000 inom jordbrukssektorn behövs det inte med nödvändighet större ekonomiska resurser , när allt kommer omkring .
man måste också göra besparingar .
men det rör sig om intellektuella resurser : man måste investera i humankapital .
det är nämligen nödvändigt att uppnå två mål , att vidmakthålla den europeiska modellen med ett allsidigt jordbruk , och detta måste ske på ett sätt som underlättar den fria världshandeln med jordbruksprodukter , vilket framför allt gynnar utvecklingsländerna .
det är inte lätt att kombinera dessa två mål , och det är inte självklart hur det skall gå till .
eventuellt finns det motsättningar mellan de båda målen , och det finns ingenting som tyder på att kommissionen har uppmärksammat dessa motsättningar och hur de skall lösas .
i fråga om den andra aspekten av agendan , herr kommissionsordförande , den som gäller sammanhållning och regional utveckling , kan vi förvisso uppvisa stora framsteg , men vi har fortfarande efterblivna områden , i synnerhet öområden , som man borde ägna större uppmärksamhet .
och i fråga om fisket finns det ingenting i ert program som antyder att det rovfiske som hotar att utrota hela fiskarter kommer att få konsekvenser i framtiden .
det behövs kanske större uppmärksamhet och mera esprit de finesse i dessa frågor .
fru talman ! jag vill inleda med att förstärka den varning som många kollegor uttryckt här om denna femårsplan .
när vi lägger fast mycket ambitiösa , långsiktiga mål får vi inte glömma nuet .
det var något som ledaren för min grupp , poettering , underströk i sitt inledande anförande .
unionen skall inte ta på sig en rad nya arbetsuppgifter utan att den centrala grundstommen finns för en framgångsrik europeisk ekonomi .
den grundstommen är uppenbarligen den inre marknaden .
hur starkt etablerad är den inre marknaden just nu ?
jag vill påminna prodi och de av hans kollegor som fortfarande är här om kommissionens egen undersökning av 3 000 europeiska företag .
nästan 40 procent av företagen i denna undersökning meddelar att de fortfarande har extra omkostnader för att göra produkter eller tjänster förenliga med nationella specifikationer .
detta är kommissionens egen undersökning .
detta är klassiska symtom på att nationella regeringar fortsätter att skapa hinder - byråkratiskt myndighetskrångel som hindrar marknadstillträde .
kommissionens program visar en störande belåtenhet över genomförandet av den inre marknaden .
vi måste fortsätta att utöva påtryckningar på alla områden genom att ta bort ytterligare hinder , öka pressen på de medlemsstater som underlåter att sätta den inre marknadens bestämmelser i kraft och naturligtvis utvidga till viktiga nya områden som finansieringstjänster .
endast med den inre marknaden som stark grundstomme kommer dagordningen för utvidgningen att kunna lyckas .
ett utvidgat europa måste byggas på unionens nuvarande starka sidor .
en inre marknad som täcker den utvidgade unionen kommer att vara en fantastisk prestation .
jag avslutar med att säga på alla mina konservativa kollegors vägnar - och vi är den näst största nationella delegationen i detta parlament - att vi lovar vårt fulla stöd till kommissionen och till prodi för att de skall lyckas med denna historiska uppgift .
fru talman , herr ordförande , kära kolleger ! vid omröstningen om er tillsättning stämde vi möte med er i dag .
det är nu som de seriösa frågorna börjar , eftersom vi i dag skall uttala oss om ert program .
när det gäller ert inlägg inför kammaren låt mig inrikta mig i mitt uttalande på det som ni kallade det nya ledningssättet . ni gör det till ett redskap för försoning med våra medborgare .
men bakom denna term &quot; nytt ledningssätt &quot; verkar helt enkelt frågan om institutionernas funktion ligga och frågan om våra offentliga myndigheters funktion , om vi är överens om att anse att europeiska unionen bör vara en offentlig myndighet .
bandet mellan unionens institutioner , medlemsstaternas befogenheter och de lokala och regionala myndigheterna , det går väl an .
men är det verkligen så vi kommer att försona medborgarna och den europeiska uppbyggnaden ?
är det verkligen så vi kommer att svara på de grundläggande frågorna som inte i så hög grad är &quot; vem gör vad &quot; utan snarare &quot; vad gör vi tillsammans &quot; ?
för det är just det som är problemet hos våra medborgare .
i ert uttalande tog ni upp de utmaningar som väntar oss , globaliseringen , utvidgningen och jag vill tillägga framtiden för vår sociala modell .
därför framhåller vi så starkt med min grupp detta förslag till stadga för det tycks oss att om vi skrev in utformningen av denna stadga om grundläggande rättigheter i vår tidsplan är det just för att vi står vid en historisk mötespunkt , och att unionen behöver omdefiniera de värden kring vilka den byggdes upp inom de aktuella gränserna , men också inför de kommande utvidgningarna som vi önskar så hett , men inte på vilka villkor som helst .
våra medborgare väntar sig mera europa av oss , men inte vilket europa som helst .
de förväntar sig inte att vi skall anpassa oss till globaliseringen , men att vi på grundval av vår sociala modell skall vara en organisationskapacitet för globaliseringen .
ur den synpunkten bör jag säga er att när ni engagerar er till förmån för en politisk union - och vi är positiva till den politiska unionen - kan detta inte göras om den inte grundas på vår sociala modell och det som utgör vår originalitet och vår kapacitet att bättre styra världens affärer .
fru talman , herr kommissionsordförande , fru kommissionär , herrar kommissionärer , värderade kolleger !
jag vill börja med ett citat : &quot; kommissionen kommer att fortsätta förberedelserna för en europeisk stadga för grundläggande rättigheter och lägga fram förslag för att genomföra ett ambitiöst program .
kommissionen kommer särskilt att föreslå att en äkta europeisk asyl- och invandringspolitik tas fram , och uttalar sig för att rättshjälpen och rättssamarbetet förstärks och att ett effektivt tillvägagångssätt utvecklas för att bekämpa varje form av brottslighet . &quot;
detta dokument är en fars i all sin korthet !
en fars därför att vi känner till och uppskattar kommissionär vitorinos arbete , och det som här läggs fram på papperet står därmed i klar motsatsställning till fakta .
ett sådant dokument är överhuvud taget inte någon basis för ett poängsystem .
det har prisats och lovats som en stor prestation , men jag håller fast vid att vi behöver en grund för ett poängsystem .
vi vill som parlament seriöst diskutera den framtida utvecklingen inom detta politiska område på grundval av ett program .
det vi förväntar oss är miniminormer i asylförfarandet , för att få snabb hjälp åt flyktingarna men också för att skapa klarhet för dem som inte befinner sig på flykt .
vi vill ha instrument för att förhindra missbruk .
vi vill ha en utveckling av invandringspolitiken i gemenskapen , som naturligtvis också inkluderar medlemsstaternas integrationsförmåga , och vi behöver en utbyggnad av exempelvis europols operativa uppgifter , för att här konkret vidta åtgärder för att bekämpa den organiserade brottsligheten .
vi befattar oss seriöst och mycket intensivt med dessa uppgifter , och vi förväntar oss samma sak från kommissionens sida , även om de bara handlar om att lägga fram dokument !
jag vill ta tillfället i akt och ta upp frågan om världshandelsorganisationen ( wto ) , ett område där viss överensstämmelse råder mellan kommissionens dokument och den socialdemokratiska gruppens ståndpunkt , något , som vi redan har hört , inte händer på andra områden .
det råder en viss överensstämmelse eftersom vi är för ett handelsutbyte på internationell nivå , men vi är för ett sådant handelsutbyte främst tack vare inrättandet av gemensamma lagar , gemensamma regler som kan reglera världshandeln kring ett och samma mål : att handeln skall främja tillväxten , och framför allt att tillväxten blir harmonisk där medborgarnas värde inte bara är något med ensamrätt för de mera dynamiska och konkurrenskraftiga regionerna i världen .
å andra sidan , vad är det för principer vi vill visa med ett sådant konstaterande ?
på världshandelsorganisationens nivå har den här regleringen och de här normerna lett till ett ökat handelsutbyte , det vill säga ökad rikedom , men när vi kontrollerar hur rikedomen har fördelats måste vi tyvärr konstatera att avståndet blir allt större mellan världens rikare länder och block och de fattigare och mera underutvecklade länderna .
därför är vi såväl berättigade som tvungna att ställa oss följande fråga : vad tjänar de nuvarande gemensamma lagarna till , de nuvarande gemensamma reglerna ?
vad tjänar de nuvarande förhandlingarna till , såsom de genomförs , och världshandelsorganisationens nuvarande verksamhet som å ena sidan ökar handelsutbytet , men samtidigt genererar skillnader och ökar avståndet mellan de rika och de fattiga länderna ?
vi sade därför att vi var positivt inställda till kommissionens strategi inför förhandlingarna i seattle och följande .
vi är framför allt för den strategiska visionen , men det krävs mod och djärvhet .
å ena sidan måste vi kräva att de sociala och miljömässiga rättigheterna samt konsumentskyddet införlivas i de nära förestående förhandlingarna .
det är dock först och främst fråga om att ha en långsiktig ambitiös och modig vision när det gäller reformen , inte bara av wto , utan också av internationella arbetsorganisationen ( ilo ) och förenta nationerna , men framför allt av de finansiella institutionerna , i första hand internationella valutafonden ( imf ) och världsbanken .
vi måste vara modiga och inte titta partiskt på globaliseringen , vi måste i stället ha mod att på ett globalt sätt se till att rikedomarna inte bara tillfaller de mera utvecklade länderna , utan alla världens regioner skall få en harmonisk tillväxt och utveckling .
fru talman ! även jag vill lovorda kommissionens initiativ att lägga fram en rapport om sina strategiska mål för de närmaste fem åren , även om jag hoppas att man har för avsikt att i senare dokument rätta till det överdrivna antalet generaliseringar och den diffusa prägeln på det dokument som vi behandlar i dag .
mot bakgrund av detta , fru talman , vill jag än en gång framföra min klagan över frånvaron av en fiskeripolitik .
det är överraskande att inte kommissionen som ett strategiskt mål för de närmaste åren beslutar om en process med en granskning av denna fråga inom gemenskapspolitiken , inför den reform som bör äga rum år 2002 .
denna granskningsprocess är , utan tvekan , en av de viktigaste händelser som kommer att påverka fiskesektorn under många år .
men det verkar den inte vara för kommissionen , som är ansvarig för att innan utgången av år 2001 inför rådet och parlamentet lägga fram en rapport om gemenskapens fiskeripolitik det senaste årtiondet , mot bakgrund av vilken rådet bör fatta lämpliga beslut om en förändring av denna .
faktum är att en granskningsprocess redan har påbörjats av många yrkesgrupper och institutioner , till exempel av europaparlamentet , som redan 1998 sammanställde och antog ett betänkande där de aktuella problemen och bristerna inom gemenskapens fiskeripolitik påvisades .
vi har flera gånger bett om en minimikalender för denna granskning , men vi har inte fått något svar .
två år minst är ingen lång tid med tanke på den besynnerliga situationen för fiskeripolitiken vad gäller bestämmelserna på den inre marknaden och på att missförhållandena måste lösas inom detta reformförfarande .
därför ber jag , fru talman , herr kommissionsordförande , att denna fråga , som är av stor betydelse för en så pass viktig sektor inom europeiska unionen , beaktas i denna strategi och i de strategiska målen för de närmaste fem åren .
fru talman ! jag skulle också vilja gratulera till kommissionsordförande prodis program .
jag välkomnar särskilt hans erkännande om att denna rättskaffens kammare har upprätthållit tillväxt : informationssamhället på en växande europeisk marknad och dessutom en enda helt fungerande valuta som skall ge oss möjligheten att verkligen främja välfärd , innovationsföretag , entreprenörsandan och - viktigast av allt - arbeten av maximalt varaktigt värde för våra europeiska medborgare .
jag har en iakttagelse , inte kritik , att redovisa beträffande kommissionsordförande prodis uttalande i morse som var ganska tandlöst om den ekonomiska politikens verkliga innehåll .
vi får inte ta någonting för givet i fråga om hur vi kan omstrukturera den europeiska ekonomin .
när allt kommer omkring , vad är social rättvisa om där inte finns full sysselsättning ?
full sysselsättning är det bästa sättet att skapa social rättvisa för v åra medborgare .
detta är den centrala fråga som vi skall inrikta oss på .
jag vill gärna framföra min uppskattning av ett eller två initiativ som kommissionen redan har lagt fram och som skall hjälpa oss : i synnerhet att kommissionär liikanen förbundit sig att föra en nytänkande kunskapsbaserad ekonomi .
ja , e-europa kommer att vara framtiden för oss och hjälpa oss att skapa ny välfärd och nya jobb .
jag välkomnar kommissionens initiativ nu och tidigare om stöd till våra små och medelstora företag , och jag skulle vilja gratulera vårt portugisiska ordförandeskap för dess initiativ att införa en stadga för småföretag .
det är viktigt och något som kan behandlas på toppmötet i lissabon .
jag välkomnar också kommissionär busquins idé om att skapa ett gemensamt forskningsområde för hela europeiska unionen .
detta är återigen ett sätt för oss att medverka till att skapa bättre möjligheter till sysselsättning och välfärd .
ni sade i er sammanfattning , kommissionsordförande prodi , att avreglering , konkurrensmöjligheter , lågt hållen inflation , innovation , vetenskap och teknik är viktiga faktorer för att den europeiska ekonomin skall bli framgångsrik och för att lyckas med att skapa nya jobb i framtiden .
jag håller verkligen med er om det , men vi kan inte ta något för givet .
det finns fortfarande mer som vi måste göra och toppmötet i lissabon skall bli en del av det .
så med dessa kommentarer vill jag gärna gratulera er till programmet och önska det all framgång .
fru talman , herr kommissionsordförande ! jag vill koncentrera mig på två punkter , som inte har nämnts i ert program .
jag har fått det intrycket att detta strategidokument från kommissionen för de närmaste fem åren skall läsas som ett vetenskapligt arbete om europeiska unionen , eller som en principförklaring .
men den ger inte intryck av någon verklig politisk strategi från kommissionens sida .
som kultur- och utbildningspolitisk talare för min grupp hade jag dessutom av just en italiensk kommissionsordförande kunnat förvänta mig mer innehåll .
på detta vis ger inte kommissionen europa någon själ !
det finns inte alls någon kultur eller utbildning i detta dokument . men det är nödvändigt att skapa ett verkligt europeiskt utbildnings- och kulturområde .
bara ett par stickord .
jag talar om att införliva kulturindustripolitik i detta utbildnings- och kulturområde ; den skapar arbetstillfällen .
jag talar om att skapa en kulturell mainstreaming på alla politiska områden , om att förstärka och förbättra den europeiska inriktningen på innehållet i utbildningen , liksom om att knyta samman utbildningspolitiken i europa . jag vill understryka det livslånga lärandet .
herr kommissionsordförande ! ni talade inte heller om det europeiska audiovisuella området , och detta i början av det nya århundradet !
dessutom konstaterar jag att informationspolitiken och kommunikationen , som bör anpassas till medborgarnas behov , inte heller nämns .
jag tror alltså att det fattas något i detta program .
ett verkligt europeiskt medborgarskap är beroende av att ett verkligt utbildnings- och kulturområde skapas och synliggörs .
principförklaringar räcker inte !
vi behöver innehåll som kontinuerligt genomförs av kommissionen på det sätt som jag tidigare förklarade , genom politiska åtgärder .
fru talman ! herr prodi , hur skulle då sammanfattningen av er politik , ert arbetsprogram och er måttstock se ut om ni var tvungen att ställa upp i direkta val ?
ni har den goda , charmanta idén att resultatet och måttstocken för er politik och för ert femårsprogram kommer att avgöra valresultatet respektive valdeltagandet vid nästa europaval .
om jag föreställer mig att jag skall presentera ert arbetsprogram för mina väljare , som jag träffar varje vecka och som jag varje vecka måste förklara det för - inte på högre politisk nivå , utan på gatan - då frågar jag mig vad jag skall säga ?
herr prodi , vad skall jag säga att det finns för nyheter i det ?
det finns ingenting nytt i ert arbetsprogram .
för fem år har ni använt 12 sidor , för ett års arbetsprogram har ni använt 18 sidor .
ger det mig några förhoppningar för år 2000 ?
nej , det gör det inte !
i ert arbetsprogram 2000 säger ni något mycket klokt .
ni säger att miljöhänsyn måste integreras i alla andra politiska områden .
har ni gjort det , herr prodi , och har ni också läst årets arbetsprogram ?
ni har nämligen inte gjort det !
ni har inte integrerat miljöpolitiken i utvidgningen , fastän det är ett av kärnproblemen i samband med utvidgningen .
ni har inte heller integrerat den i den ekonomiska politiken , konkurrensen eller den inre marknaden .
ni har inte gjort det någonstans .
ni har sammanfogat enskilda sättstycken , men ni har inte skapat någon helhet .
ni sade tidigare i ert tal att en sådan katastrof som den som skett i donau måste ge anledning till ett katastrofprogram - nej , herr prodi , vi måste äntligen börja genomföra lagstiftningen och även se till att vi kan kontrollera lagstiftningen .
ni skriver i ert femårsprogram att människorna i europeiska unionen med all rätt förväntar sig bättre livsmedelsstandarder och bättre livsmedelslagstiftning .
herr prodi , ni vet inte vad ni talar om !
europeiska unionens livsmedelslagstiftning är den mest ambitiösa i världen !
det som saknas , är att den skall genomföras och kontrolleras i medlemsländerna .
ta äntligen er uppgift på allvar att som ordförande för kommissionen ta medlemsstaterna i öronen och tvinga dem att göra sin plikt och genomföra sina uppgifter !
de skall inte alltid bara ägna sig åt sina fritidssysselsättningar , utan utföra det dagliga normala arbetet .
det förväntar vi oss av er under de närmaste fem åren !
fru talman , herr kommissionsordförande , mina damer och herrar ! ni gör det inte enkelt för mig som ordförande för fiskeriutskottet , herr prodi .
jag ser mig tvungen att offentligt här i dag kritisera fiskets frånvaro i det program som ni har lagt fram .
de närmaste fem åren kommer prodis kommission - detta tillkännager ni högtidligt i den första av era slutsatser - att genomgå stora förändringar .
jag hoppas att de förändringar som ni tillkännager inte innebär en ännu större diskriminering av fisket , att döma av den väldiga och totala tystnad som frågan omges av i ert program .
inte en rad , inte ett ord angående fisket eller den gemensamma fiskeripolitiken .
jag begär inga detaljer eller konkretiseringar , men jag anser att ett omnämnande vore på sin plats .
hur är det möjligt att en gemensam - jag upprepar , gemensam - politik med en sådan ekonomisk , social och regional genomslagskraft - och som påverkar europas ekonomiska och sociala sammanhållning , har blivit bortglömd ?
ännu värre , om möjligt med tanke på att kommissionen , herr prodi , - så som påpekades - skall genomföra granskningen eller reformen av den aktuella gemensamma fiskeripolitiken , som den är ålagd att göra år 2002 .
kommer inte kommissionen heller att göra något - åtminstone tillkännages inget sådant - år 2000 åt denna reform ?
vilket är då budskapet till europas fiskare , till deras familjer och till fiskeriindustrin , såväl själva fisket som dess bearbetande och saluförande grenar , och till närbesläktade eller stödjande industrier som är beroende av fisket i så och så många europeiska hamnar i så och så många europeiska regioner , många av dem för övrigt i ytterområden , som med all rätt kräver att man fokuserar uppmärksamheten på detta problem ?
ni hänvisar inför de närmaste åren tydligt till den gemensamma jordbrukspolitiken , men ni säger inget om den gemensamma fiskeripolitiken vad gäller den dubbla anpassning som måste ske av den inre marknaden för att det inte skall finnas några undantag - något som också har påpekats här - i ett globalt sammanhang , i denna globalisering .
parlamentet har uttalat sig på den första punkten och kommer också att göra det på den andra .
jag ber er därför , herr prodi , att ni tar upp detta i ert svar i dag .
vår parlamentsgrupp kommer att lägga fram ett ändringsförslag i den frågan och jag skulle vilja att ni gav oss ett positivt besked .
herr kommissionsordförande ! det här är ett historiskt ögonblick för parlamentet , ett femårsprogram efter kommissionens kris .
jag skulle för den socialdemokratiska gruppens räkning vilja koncentrera mig på punkten angående inre reformer .
vi stöder gärna programmet så som det nu lagts fram i en samrådsakt och som även återkommer i vice ordförande kinnocks program för kommissionens räkning .
vi tycker det är mycket viktigt att vi , när det gäller ekonomisk kontroll , personalpolitik och kortare byråkrati , ser fram emot snabba beslut och en effektivare byråkrati , till medborgarnas tjänst .
samtidigt inser vi att det är ett enormt stort program och att under de kommande årens ombyggnad så måste samtidigt butiksförsäljningen fortsätta med konkreta resultat .
på samma sätt som kvinnorna i nederländerna plötsligt upptäckte att de kunde hänvisa till den europeiska lagstiftningen för att de låg för långt efter med avseende på den sociala tryggheten , gäller i dag också samma sak för flera andra medborgare .
demokrati , öppenhet , insyn och tydlighet hör alltid ihop med resultat , medborgare uppskattar resultat och det är på dessa som kommissionen bedöms .
det är precis som kollega swoboda och även andra kolleger här redan sagt : rädslan för modernisering , globaliseringen , den enskilda personen som förlorar sin egen trygghet och säkerhet .
det kan förebyggas med hjälp av den europeiska sociala modellen och om resultat uppnås på alla de här konkreta områdena .
mitt innerliga yrkande för stöd till den inre reformen hör alltså lika mycket ihop med konkreta resultat på det sociala området , så att medborgaren känner igen sig , här i europa och även där utanför .
den medborgaren , en femtedel av världsbefolkningen , har fortfarande inte tillgång till grundläggande sociala möjligheter som till exempel undervisning och hälsovård .
det är dessa som vi verkligen måste visa solidaritet med .
fru talman , ärade kommissionsordförande , ärade kollegor ! jag har läst och återigen läst kommissionens dokument om de strategiska målen för mandatperioden .
det gläder mig att vi har diskuterat det i parlamentet , jag noterar löftena och jag noterar det som utlämnats .
kommissionen nämner bara helt apropå den ekonomiska och sociala sammanhållningen , solidariteten mellan medlemsstaterna och europeiska unionens regionala politik , och detta samtidigt som man tar upp utvidgningsfrågan .
kan det vara så att målet skall anses vara uppnått med en mindre skillnad mellan tillväxtnivå och det påföljande stödet för den faktiska konvergensen ?
med all säkerhet inte !
under tiden menar man mycket riktigt att europa måste omvärdera rollen som solidarisk partner till u-länderna samt koncentrera sig i kampen mot fattigdomen .
vad stort sker , det sker tyst .
kommissionens sätt att inte ta upp sammanhållningen är för mig allvarligt .
man förringar en princip i fördragen - den ekonomiska och sociala principen - som skall genomsyra all politik och alla åtgärder vidtagna av de europeiska institutionerna , man verkar vara ovetande om att många europeiska regioner är kraftigt underutvecklade , man glömmer att utvidgningen rättfärdigas av ett gott omdöme i den regionala politiken .
utan verklig konvergens är sammanhållningen inom europeiska unionen i fara .
kom ihåg den sjätte periodiska rapporten om tillståndet för europeiska unionens regioner , som kommissionen är ansvarig för .
med en genomsnittlig tillväxtnivå på 100 konstaterar man att de tio regioner som anses vara de &quot; starkaste &quot; i genomsnitt ligger på 158 , och de tio &quot; svagaste &quot; stannar på 50 .
dra era egna slutsatser .
50 : just den tillväxtnivå som min region , azorerna , hamnade på - en av dem som i fördragen definieras som en ultraperifer region .
jag väntar på kommissionens betänkande om ultraperifera regioner som rådet fastslog skulle utarbetas till december 1999 .
jag slutar med att på nytt påtala min övertygelse : utan ekonomisk och social sammanhållning kommer ingen sammanhållning alls att uppnås , bara upplösning .
fru talman , herr ordförande !
vi och den europeiska allmänheten behöver en stark kommission , för enligt fördragen och också folkets vilja är kommissionen motorn i den europeiska uppbyggnaden , den sisyfosklippa som vi tillsammans måste bära upp till toppen igen efter varje utvidgning .
således , en stark kommission men som stöder sig på parlamentet , och parlamentet är således er allierade , men det är en besvärlig allierad vars meddelanden bör avlyssnas och jag skulle vilja lämna några meddelanden i detta korta inlägg .
för det första , herr ordförande tror jag att även om era båda föregångare huvudsakligen ägnade sig åt att utveckla en inre marknad och inrätta en gemensam valuta är det huvudsakligen er sak att utveckla det medborgarvärde som står i centrum för den europeiska uppbyggnaden .
ni får nämligen inte låta er distraheras enbart av utvidgningsärendet , hur viktigt det än är .
ni måste gå längre i riktning mot en försoning av medborgarna med europa och i synnerhet de medborgare som är offer för ekonomiska , sociala och otvivelaktigt på sikt tekniska brytningar .
främjandet av vetenskaplig utveckling , även främjandet av nya tekniker och allas tillgång till dessa tekniker kommer inte att säkras av marknaden och av konkurrensen , inte mer än att marknaden och konkurrensen kommer att säkra den sociala närheten och effektiviteten när det gäller de stora kollektiva tjänsterna , hälsa , utbildning , transporter , kommunikationer , vatten och jag vet inte vad .
ert åtgärdsprogram och era målsättningar är diskreta och rentav helt tysta när det gäller konsolideringen och finansieringen av de stora offentliga tjänsterna och tjänster av allmänt intresse .
det finns en absolut prioritering , herr ordförande , om ni vill försona europa med medborgarna : att se till att de hellre väljer europa än jörg haider .
fru talman ! kommissionen gjorde rätt när den gjorde livsmedelssäkerhet till en av de viktigaste frågorna .
den nyligen inträffade dioxinskräckhistorien i belgien , den tidigare bse-krisen i storbritannien och den pågående kontroversen om hur farliga genetiskt modifierade livsmedel är har alla bidragit till att konsumenterna litar mindre på att den mat de äter är ofarlig .
om kommissionen verkligen kan återställa förtroendet för livsmedelsproduktionskedjan kommer den samtidigt att återskapa förtroendet för europeiska unionens institutioner och visa deras förmåga att skydda eu-medborgarnas rättigheter .
jag välkomnar därför det faktum att frågan om livsmedelssäkerhet , folkhälsa och konsumentförtroende understryks markant i kommissionens arbetsprogram för år 2000 .
jag blev dock besviken över hur förslaget om inrättandet av en europeisk livsmedelsmyndighet är utformad i den senaste vitboken .
i dess nuvarande form är det som föreslås mer som ett rådgivande organ till kommissionen snarare än ett självständigt organ som skulle ha beslutande och lagstiftande befogenheter mer likt dem hos den amerikanska livsmedelsmyndigheten : food and drug administration , vilken redan har skapat trovärdighet på detta speciella område .
vidare måste man i det framtida lagstiftningsarbetet ta itu med arbetsmetoden för samspelet mellan den europeiska livsmedelsmyndigheten och myndigheterna i nationella medlemsstater , exempelvis myndigheten för livsmedelskontroll i irland .
detta organ , exempelvis , utför tillsammans med det nyligen inrättade gränskontrollorganet i irland för livsmedelssäkerhet redan ett bra arbete .
det skulle vara tragiskt om deras ansträngningar skulle undergrävas på grund av brister i eu : s lagstiftning .
jag fruktar att sådana brister i eu : s lagstiftning kan leda till revirstrider mellan nationella organ och eu-organ , som borde arbeta tillsammans i stället för att mot varandra .
det är något som vi måste bevaka .
fru talman ! ordförande prodis presentation i dag var nödvändigtvis en ganska brett svepande historia .
vi kommer att titta efter enskilda detaljer år för år , till exempel i det sociala åtgärdsprogrammet som skall läggas fram i år .
vi skall också granska detta från perspektivet social- och sysselsättningspolitik och genomföra en rad kontroller .
vi skall granska i vilken omfattning vi kan skapa en liksidig triangelformad politik där man kombinerar ekonomisk politik , sysselsättningspolitik och socialpolitik .
för ögonblicket ligger socialpolitiken långt bakom politikområdena ekonomi och sysselsättning .
inom ramen för sysselsättningsstrategin skall vi sträva efter att fördjupa och bredda strategin efter översynen under det portugisiska ordförandeskapet och inom den ram som förslagits av det portugisiska ordförandeskapet .
inom ramen för den sociala dimensionen skall vi sträva efter att fördjupa den inre marknaden med en social aspekt .
strömmen av sammanslagningar , fusioner och överlåtelser som vi upplever när marknaden får allt större intresse innebär att vi måste göra något för att aktualisera den mall för de informations- och samrådsdirektiv som vi antagit tidigare ; men vi måste också komplettera dem med det nya generella regelverket för information och samråd och uppdatera företagsrådsdirektivet .
vi behöver även en uppförandekod för bolag för att se till att företag i själva verket arbetar i partnerskap med sina anställda i förändringsarbetet .
det är ett framgångsrikt sätt att hantera förändring och jag hoppas kommissionen kommer att se till att det genomförs .
slutligen , med uppdykandet och återuppvaknandet av rätten till främlingsfientlighet inom europeiska unionen hoppas jag att våra institutioner tillsammans kommer att göra sitt yttersta för att ge artikel 6 verkligt innehåll genom att tillämpa artikel 13 för att bekämpa diskriminering och artikel 137 för att bekämpa uteslutning .
vi måste snarast börja arbeta med den dagordningen nu .
förhoppningarna , ordförande prodi , är bra men vi vill att dessa förhoppningar skall paras med åtgärder .
fru talman ! jag hoppas att det är ett gott tecken att jag avslutningsvis får påpeka ytterligare en sak !
herr prodi , i era reformsträvanden är ni särskilt intresserad av att förverkliga en framtidsorienterad sysselsättningspolitik över hela europa .
men för just den ekonomiska sektor som jag företräder , fiskerisektorn , betyder detta förändringar .
vi måste överge de planekonomiska subventionerna och komma fram till en liberal politik , som främjar det egna ansvaret .
vi måste sänka skyddstullarna för att garantera att företagen inom tillverkningsindustrin tas i anspråk effektivt .
så handlar det slutligen om det europeiska näringslivets konkurrenskraft på världsmarknaden och om tusentals arbetstillfällen inom tillverkningsindustri och havsfiske .
men jag behöver säkert inte påminna er om betydelsen av en näringsgren som inte bara är en nationalekonomisk faktor , utan också en samhällsfaktor , som inte bara berör tyskland , utan gränsövergripande berör alla kustregioner i europa .
dessutom är denna näringsgren en av de få sektorer som fullt ut har integrerat europeiskt besluts- och handlingsansvar . därför förväntar vi också här att vi får medbeslutanderätt .
det rekommenderas nu enhälligt .
men revideringen av fiskeripolitiken är fastställd till att äga rum om några månader , dvs. i början av år 2000 .
då är det verkligen störande att denna näringsgren alls inte nämns i föreliggande dokument .
jag hoppas att det här handlar om ett missförstånd !
jag ber , herr prodi , att stå för vad ni sagt , och genomföra det !
fru talman ! många av talarna från socialistgruppen har redan identifierat viktiga områden där det finns brister i kommissionens uttalande .
vi har dock uttryckt att detta är ett nyskapande och mycket välkommet initiativ av kommissionen .
ett område som jag vill inrikta mig på , förutom dem som redan nämnts , är kulturell mångfald i europa .
i inledningen till detta uttalande tillstås i avsnittet om livskvalitet att detta är viktigt .
men det finns inget i uttalandet som visar att kommissionen avser att vidta några åtgärder för att hantera frågan om kulturell mångfald .
om vi skall kunna garantera att vi besegrar dem som sprider rädsla ibland oss - dem som strävar efter makt med stöd av oroliga medborgare - då måste vi allvarligt ta itu med frågan om hur vi kan leva tillsammans och hur vi kan undanröja de negativa stereotyper som vi har om varandra , både inom den nuvarande europeiska unionen och bland dem som försöker ansluta sig och rent av bland dem i andra delar av europa och världen som vill komma hit och bo och arbeta i europa .
om vi inte tar itu med dessa frågor , om vi inte kan undanröja dessa negativa stereotypa uppfattningar , om vi inte använder det som är bäst från våra olika kulturer och språk och skyddar och utökar det och ser till att vi menar allvar med att ha ett mångfaldigt europa , kommer vi att misslyckas .
de som just nu är i blickpunkten i europa grundat på rädsla skall vinna slaget .
jag är allvarligt oroad att om kommissionen inte inser att detta är en viktig aspekt på hur vi skall skapa ett samhörande europa kommer vi att göra framsteg på det ekonomiska området och på sysselsättningsområdet och även inom utrikes- och säkerhetspolitik men våra medborgare kommer fortfarande att vara ängsliga därför att de kommer att vara rädda för det okända och rädda för dem som de inte förstår .
om vi inte vidtar åtgärder för att hantera detta kommer vi till sist att misslyckas .
kära kollega , jag tackar er .
innan jag på nytt ger ordet till kommissionens ordförande vill jag meddela er att jag i enlighet med artikel 37 har fått sju resolutionsförslag till sammanfattning av debatten .
välkomsthälsning
herr talman ! även jag vill ta upp en ordningsfråga .
finns det några regler eller förordningar som reglerar demonstrationer inom parlamentets byggnad , utanför dörrarna till kammaren , för att säkerställa att ledamöter kan komma in i denna kammare för att fullgöra sina uppdrag ?
om det finns sådana regler vem ansvarar för att de efterlevs och vad gör de för att uppfylla det ansvaret ?
herr talman ! jag skulle vilja ta upp frågan om assistentstadga igen , som vi alltid har prioriterat , och informera er om att vi - den italienska delegationen i gruppen - på gruppens ordförande barón crespos uppmaning har deponerat de kontrakt vi har upprättat med assistenterna hos kvestorerna .
jag tycker att det är en konkret gest för att komma till en lösning på detta problem .
därför skulle jag vilja uppmana parlamentets presidium att överväga om det inte vore lämpligt att presidiet uppmanade alla ledamöterna att göra detsamma .
herr talman ! låt mig först och främst säga att jag helt stöder kravet på en stadga för assistenter .
i går när jag anlände till parlamentet fick jag en skrivelse om en föreslagen demonstration av assistenterna utanför parlamentets dörrar .
som alla kollegor känner till - och många av er har kontaktat mig under de senaste sex månaderna - bedöms alla utställningar och liknande arrangemang först av parlamentets comartkommitté ( comité des arts - konstkommittén ) .
för att ge ett ej omtvistat exempel : inga kommersiella utställningar får hållas här i parlamentet av uppenbara skäl .
efter att jag mottog ett brev i går informerade jag omedelbart assistenterna att vi skulle föreslå att de fick hålla ett möte eller demonstration , förmodligen inom en snar framtid och eventuellt under nästa månad .
men alla sådana arrangemang måste genomföras på ett sätt som inte stör parlamentets reguljära verksamhet .
jag undertecknade ett brev i går eftermiddag vid parlamentspresidiets sammanträde i vilket assistenterna informerades om detta .
men jag har också hört att de informerades muntligen om detta beslut av gruppordförandekommittén i torsdag , så de var helt medvetna om beslutet .
problemet är inte att de talar om för oss hur de känner , det är inga problem med ett eventuellt möte under parlamentets nästa delsession .
men det blev ett missförstånd då de mottog ett brev från en annan person som de ansåg gav dem tillstånd .
alla utställningar blir emellertid först bedömda av den så kallade comartkommittén .
som ni vet har vi många utställningar runt om i parlamentsbyggnaden om olika länder eller om vad som helst .
detta är inte ett försök att vare sig censurera eller gå emot den mycket reella och befogade principen att vi bör ha en stadga för assistenter .
tack för det , ledamot banotti .
ert inlägg borde kunna klargöra olika frågor som har tagits upp .
vi skall nu genomföra omröstningen.1
herr talman ! jag talar som företrädare för den spanska delegationen av europeiska folkpartiets grupp ( kristdemokrater ) och europademokrater , för delegationen av det spanska folkpartiet , beträffande terrón i cusís resolution om området med frihet , säkerhet och rättvisa .
faktum är att vi inte i alla omröstningar har följt direktiven från europeiska folkpartiets grupp , och vi har röstat för terrón i cusís resolution som på det hela taget är en utmärkt resolution .
däremot röstade vi emot punkterna 2 och 6 , för vi anser att de är oriktiga juridiskt sett .
i stället har vi röstat för skäl j som ligger i linje som det jag själv , som föredragande av yttrandet , har föreslagit utskottet för medborgerliga fri- och rättigheter samt rättsliga och inrikesfrågor inför regeringskonferensen .
vi har likaså röstat för punkt 13 .
en ändamålsenlig stadga och fri rörlighet och etablering för tredje land är något som det spanska folkpartiet länge har försvarat .
av liknande skäl har vi röstat för punkt 14 där , i och med det muntliga ändringsförslaget en viss , högst berättigad oro för problem med subsidiariteten har beaktats , och där både vad gäller de politiska rättigheterna , inte längre rösterna i kommunvalen , utan de politiska rättigheterna i generella termer , ingår i medlemsstaternas suveränitet .
i och med det muntliga ändringsförslaget tyckte vi att vi kunde rösta för detta och det har vi också gjort .
( da ) de danska socialdemokratiska ledamöterna av europaparlamentet har valt att rösta för resolutionsförslaget , men betonar samtidigt att vissa områden strider mot det undantag som danmark har på det rättsliga området - ett undantag som den danska delegationen i pse-gruppen naturligtvis vill respektera .
. ( fr ) detta betänkande , som jag inte har röstat för , handlar i mindre grad om mänskliga rättigheter än om &quot; gemenskapsinförlivande &quot; , i själva verket konsolideringen av fortet europa .
de &quot; framsteg &quot; från 1999 som tas upp i betänkandet är bara framsteg i förhållande till dublinkonventionerna och schengenavtalen , och ännu en handlingsplan från tammerfors , som inskränker invandrarnas rättigheter .
för i förhållande till mänskliga rättigheter är det en tillbakagång .
europa fortsätter att avvisa personer till länder som anses farliga av fn : s flyktingkommissariat medan en del länder i central- och östeuropa som är eu-kandidater tar emot zigenarflyktingar som i mängd avvisats från belgien .
albaner från kosovo och serbiska desertörer förvägras flyktingstatus medan pinochet i lugn och ro klarar sig undan sin process .
schengenkonventionens europa jagar avgjort lättare förföljda från söder än diktatorer , samtidigt som fn anser att vi kommer att behöva 159 miljoner invandrare för att behålla den demografiska balansen från och med nu till år 2025 .
europa bör legalisera alla personer som är utan uppehållstillstånd , ge dem asylrätt och rösträtt till alla val och sedan kan vi i kammaren tala om ett område för frihet och rättvisa .
betänkande ( a5-0026 / 2000 ) av mccarthy
herr talman ! jag vill börja med att påpeka att jag som borgmästare i bilbao på nittiotalet fick tillfälle att lägga fram ett av de första urbana pilotprojekt som kommissionen skulle ge anslag till .
våra erfarenheter i bilbao av detta pilotprojekt har lett fram till fyra slutsatser : den första är att europa måste behålla en urban politik och , i stället för att minska resurserna från 900 miljoner euro under föregående femårsperiod till 700 för innevarande femårsperiod , bör öka finansieringen av programmet , till exempel - så som vi i gruppen de gröna / europeiska fria alliansen har föreslagit - genom att i urban-projekten åter investera den del av strukturfonderna som varje medlemsstat inte har förbrukat inom fastställt datum .
för det andra bör insatserna , när det är dags att besluta vilka områden man bör ge anslag till , koncentreras till projekt med en genomgripande verkan .
spridda åtgärder är inte effektiva .
man måste välja , och prioritera de värsta och mest överhängande fallen , till förmån för de fasta målen i sin helhet , det vill säga för de sociala , ekonomiska och miljömässiga aspekterna med en demokratisk förvaltning , liksom förhållandet mellan dem .
för det tredje bör man ta hänsyn till den synergism som ger upphov till andra gemenskapsprogram , liksom möjligheterna till en hållbar utveckling inom den miljö eller det område som avses .
slutligen måste man lita på de instanser som finns närmast medborgarna , nämligen kommunerna och de lokala organen och stödja dessa .
det är främst där man känner till de sociala behoven , där man är starkast engagerad i problemen och dessutom där man kan föreslå projekt och genomdriva dem på ett effektivt sätt utan att belasta dem med byråkrati och uppnå de bästa resultaten .
slutligen , av våra fyra ändringsförslag i dagens omröstning har två antagits medan de övriga två förkastades .
det tvingar oss att avstå i den slutgiltiga omröstningen , för vi inser inte varför inte miljöaspekten beaktas när det att dags att fatta beslut om vilka projekt som skall finansieras , och vi begriper inte varför man inte godtar att varje medlemsstat kan avsätta den del av strukturfonderna till urban-projekten som de inte har förbrukat i enlighet med gemenskapsprogrammen .
herr talman ! jag skulle vilja påminna om att vi har haft många diskussioner i utskottet för regionalpolitik , transport och turism om urban-initiativet .
många idéer har framförts . jag skulle också vilja påminna om att det trots allt var det minsta gemenskapsinitiativet som fanns och att vi följaktligen hade föreslagit att anslaget skulle ökas genom ett ändringsförslag , som förkastades .
vi beklagar detta eftersom det nämligen fanns kvar pengar från strukturfonderna i en del länder och dessa pengar skulle verkligen ha kunnat stödja pilotprojekt , eftersom urban-projekten , vill jag påminna om , just är pilotprojekt som gör det möjligt att genomföra en verklig politik för städerna .
jag skulle också här vilja uppmärksamma kommissionen på sammanhållningen mellan de olika politikområden som genomförts och jag skulle också vilja att kommissionen gör en sammanhållning av urban-projekten med de framtida projekten från den budgetpost som kallas &quot; hållbar stadspolitik &quot; .
jag skulle slutligen också vilja påminna om att vi i dag fortfarande inte har någon europeisk politik för städerna i europeiska unionen och jag vill klargöra att denna punkt , kanske , skulle kunna utvidgas inom ramen för omorganisationen och regeringskonferensen så att europeiska unionen äntligen också får en verklig politik för städer .
herr talman ! jag skulle vilja påpeka att jag röstade för detta betänkande om hållbar stadsutveckling , vid namn urban .
liksom alla de andra gemenskapsinitiativen är det någonting mycket positivt .
europa visar sig närvarande just i det ögonblick när man gör någonting för alla europeiska medborgare och inte bara för en enskild stads utveckling , vilken det vara må .
med urban vill man hitta lösningar på städernas förfall , och detta är någonting som intresserar de äldre mycket och som därmed intresserar pensionärspartiet mycket .
det finns ingen som har det sämre än en äldre människa i staden .
jag hoppas att detta gemenskapsinitiativ kommer att bli ett föredöme för hur man löser problemet med äldre i städerna .
( da ) vänsterns fem ledamöter av europaparlamentet har valt att stödja leader + , equal-initiativet och interreg , men inte urban .
vid en kommande granskning av dessa program bör eu : s insats koncentreras på gränsöverskridande uppgifter och anpassas till en utvidgning av eu .
vi har röstat för betänkandet om meddelandet från kommissionen om fastställande av riktlinjer för ett gemenskapsinitiativ för ekonomisk och social förnyelse av städer och förorter som befinner sig på tillbakagång för att främja en hållbar stadsutveckling ( urban ) .
i grunden är vi emot denna typ av program och strukturfonder , men eftersom omröstningen endast behandlar hur - och inte om - dessa resurser skall användas , har vi endast tagit ställning till innehållet och anser allmänt att förslaget om förnyelse av städer och förorter som befinner sig på tillbakagång innehåller förnuftiga slutsatser samt goda förslag och kriterier för projekten .
. ( fr ) i betänkandet räknas allmänna begrepp upp rörande vad som kallas en strategi för urban förnyelse av stadskärnor och förorter som drabbats av den kapitalistiska ekonomins kris och dess konsekvenser : ökad arbetslöshet , utestängning och ungdomsbrottslighet .
i betänkandet understryks att för att säkra en hållbar utveckling i städerna , gäller det att genomföra en urban politik som inte åsidosätter de främsta offren för den ekonomiska krisen : arbetslösa , invandrare , flyktingar , kvinnor och utestängda .
men det sägs ingenting om skälen och de ansvariga till krisen .
i betänkandet är det bara i bästa fall fråga om att rätta till vissa aspekter och efterverkningar av den .
och dessutom med chockerande neddragna medel , eftersom enligt betänkandet själv är anslagen som tilldelats programmet urban ii för perioden 2000-2006 omkring 30 procent lägre än anslagen från den föregående perioden , som redan var låga ( 900 miljoner euro ) trots att det handlar om ett femtiotal projekt i hela europa , vilket är obetydligt , när det är strängt taget samtliga storstadsförorter i vår världsdel och rentav stadskärnor som drabbas .
därför röstar vi regelbundet för de konkreta åtgärder som anmälts för att hjälpa de minst gynnade sociala kategorierna , men vi avstår i fråga om själva betänkandet genom att ange att det härrör från fromma önskningar som finansierats med rabatt .
( fr ) fru föredragande , mina kära kolleger ! jag måste säga att jag är mycket nöjd med att gemenskapsinitiativet urban fortsätter , ett initiativ som siktar till att stödja den sociala och ekonomiska omvandlingen i städer och förorter i kris , detta för att främja en hållbar utveckling i städerna .
med omkring 80 procent av den europeiska befolkningen boende i stadsmiljö är städerna i centrum av den ekonomiska , sociala och kulturella utvecklingen i europa .
samtidigt är de sociala och ekonomiska problem som det europeiska samhället brottas med mer markanta i städerna .
många europeiska städer har nämligen en intern regional brytning : samexistensen , i städerna , av kvarter där man bedriver verksamheter med högt mervärde och där höginkomsttagare är bosatta och av kvarter , som markeras av låga inkomster , hög arbetslöshet , medelmåttiga och överbefolkade bostäder och ett starkt beroende av socialstöd .
koncentrationen av sociala och ekonomiska problem till vissa stadsområden kräver en målinriktad intervention som tar hänsyn till problemens komplexitet .
därför har europaparlamentet krävt och lyckats uppnå en förlängning av gemenskapsinitiativet urban i reformen av strukturfonderna .
urbans framgång under programplaneringsperioden 1994-1999 är obestridlig .
resultatet är påtagligt när det gäller förbättring av livskvaliteten i de målinriktade områdena .
detta gemenskapsinitiativ främjade utvecklingen av goda metoder inom de ekonomiska , sociala och miljömässiga sektorerna .
det hade dessutom fördelen att stärka rollen för de lokala myndigheternas , icke-regeringssektorns och de lokala myndigheternas roll och främja nya partnerskapsformer på området förförnyelse av städer .
med det nya initiativet skall vi fortsätta att försöka nå dessa mål genom att stärka dem samtidigt som vi särskilt tar hänsyn till främjandet av lika möjligheter för män och kvinnor och integrationen av kategorier av människor som är socialt marginaliserade och missgynnade .
vi kan således glädja oss åt att det antagits .
man måste emellertid medge att på det finansiella planet kan vi inte utropa segern !
det avsatta finansiella totalanslaget är nämligen inte på långa vägar i nivå med det som står på spel .
anslagsbeloppet var 900 miljoner euro för perioden 1994-1999 och det är 700 miljoner euro för perioden 2000-2006 , det vill säga en minskning med 30 procent !
denna minskning av finansmedlen har lett till en minskning av antalet program inom ramen för det nya urban-initiativet .
det valda taket tycks vara för lågt . det har satts till femtio projekt .
det bör således ökas för att regionala och lokala faktorer skall beaktas samtidigt som de finansiella anslagen avsedda för medlemsstaterna behålls .
mot bakgrund av denna koncentration på ett antal begränsade projekt spelar kanske offentliggörande och spridning av resultaten från det nya gemenskapsinitiativet urban en viktig roll för att få en ökningseffekt .
. ( fr ) betänkandet mccarthy om gemenskapsinitiativet urban ger oss tillfälle att diskutera om det är lämpligt att gemenskapen ingriper på stadsområdet .
situationen i vissa stadsområden är alarmerande och den sociala nöden visar sig i form av arbetslöshet , fattigdom och kriminalitet .
narkotikahandeln i synnerhet underhåller osäkerhet och småbrottslighet .
strukturfondernas effektivitet är tvivelaktig inför sådana sociala utmaningar .
subsidiariteten borde leda till att vi erkänner att staten i utövandet av sina regeringsfunktioner och de lokala myndigheterna är mest lämpade för att ingripa på rätt sätt , staten genom att trygga den allmänna säkerheten och de lokala myndigheterna genom att hjälpa människor i svårigheter .
även om man kan glädja sig åt viljan att skapa ett system för utbyte om lyckade företag , kan man inte ställa de specifika problemen för varje stadsområde på samma plan .
gemenskapsinitiativet urban ingår i europeiska unionens vilja att införliva stadspolitiken i gemenskapen .
det skulle vara mera relevant om europeiska unionen inriktade sina finansiella ansträngningar på redan befintliga europeiska politikområden .
en del grupper och personer passar självklart på tillfället att ge sig in på ett nytt budgetöverbud , ett överbud som är speciellt illa valt vid en tidpunkt då staternas budget tvingas till en allvarlig avmagringskur på grund av emu : s konvergenskriterier .
mccarthy föreslår således en ökning av de avsatta anslagen till urban och främjande av detta gemenskapsinitiativ genom en dyrbar kommunikationskampanj som kommer att användas till att berömma det federala europas goda gärningar .
måste man påminna om att en utgifts effektivitet inte mäts i storleken på de anslag som tilldelas projektet ?
däremot anser mottagarna av alltför många och höga subventioner att dessa på sikt kan tas för givna .
målsättningen bör inte vara att stödja medborgarna utan att få dem att ta ansvar .
i betänkandet betonas slutligen starkt åtgärder till förmån för etniska och sociologiska minoritetsgrupper .
vi kan bara förkasta en minoritetspolitik som ofrånkomligen är farlig för den sociala sammanhållningen .
å ena sidan , uppmuntras genom denna politik till integration av invandrare där det skulle vara nödvändigt att främja deras assimilering med mottagarlandets kultur för att undvika att etniska getton uppstår som blir en explosionsrisk i staden .
å andra sidan , laborerar den med principen om positiv diskriminering , en politiskt korrekt illusion och minst lika skadlig , såsom den amerikanska presidenten har visat .
på grund av dessa orsaker kunde den franska delegationen i uen-gruppen inte godkänna betänkandet mccarthy .
betänkande ( a5-0028 / 2000 ) av decourrière
herr talman ! programmet interreg ligger oss särskilt varmt om hjärtat .
jag gläder mig liksom många av mina kolleger åt att parlamentet har kunnat behålla detta interreg-initiativ .
eftersom jag själv bor i området sarre-lorraine-luxemburg i södra belgien vet jag att det är där europa skapas , där vi lever med europa dagligen och medborgarna faktiskt ser till att den europeiska uppbyggnaden lever fullt ut .
dessa förslag bör verkligen beaktas och hållbar utveckling bör redan införlivas i dem .
varför påpekar jag det ?
helt enkelt för att de förslag som nu läggs fram fortfarande alltför ofta är miljöförstörande , på det sätt som de läggs fram .
att godkänna nya vägar , till exempel , det är att godkänna nya skadliga faktorer i europeiska unionen och det går helt emot den politik , som vi föreslår , i fråga om kamp mot gasutsläpp med växthuseffekt , till exempel .
jag ber också att kommissionen inom ramen för de projekt som läggs fram skall vaka över att miljöpelaren i europeiska unionens politik införlivas i dessa projekt och att målet att minska , till exempel , koldioxiden skall kunna vara ett pilotmervärde i de föreslagna projekten .
jag tänker här särskilt på vissa infrastrukturer som håller på att genomföras .
man vet att vissa medlemsstater fortfarande tvekar , till exempel , mellan järnväg och landsväg för genomfarter i känsliga områden såsom pyrenéerna - jag tänker på aspe-dalen .
men jag tänker också på min region där min medlemsstat fortfarande tvekar mellan att bygga järnväg och en andra motorväg , a32 .
sålunda också här ber jag således kommissionen att vara särskilt uppmärksam så att det blir en verklig sammanhållning mellan de olika politikområdena , i synnerhet i de framlagda interreg-programmen .
herr talman ! jag röstade för decourrières betänkande om gemenskapsinitiativet interreg , framför allt på grund av det svar kommissionär barnier gav några ledamöter som begärde att man i detta program skulle bry sig mer om de gränsregioner som har havsgränser .
detta gjorde jag inte bara för att jag är född i en kuststad , genua , utan framför allt för att även de gränser som utgörs av vatten är gränser .
dessa gränser vetter mot afrikas länder och mellanöstern : vi måste ta större hänsyn till det faktum att det är viktigt att utveckla också kustregionerna i alla delar av europa .
. ( fr ) i min egenskap av ledamot av europaparlamentet från ett gränsområde emotser jag med stort intresse det tredje interreg-initiativet .
vi kan aldrig tillräckligt påminna om de svårigheter som fanns förr i tiden i de områden vid gränserna , på land eller till havs , som hade delats ekonomiskt , socialt och kulturellt .
på grund av närvaron av gränser omvandlades de till yttersta randområden i de stater där de ingick , vilket alltför ofta ledde till att de statliga myndigheterna åsidosatte dessa områden inom ramen för den nationella politiken .
därför infördes gemenskapsinitiativet interreg från och med 1990 .
syftet med programmet var att uppmuntra till gränsöverskridande , transnationellt och interregionalt samarbete samt en balanserad utveckling av gemenskapens område för att stärka den ekonomiska och sociala sammanhållningen i unionen .
interreg syftar huvudsakligen till att finansiera gemensamma metoder för utveckling av små och medelstora företag , yrkesutbildning , grundutbildning , kulturellt utbyte , hälsofrågor , miljöskydd och miljöförbättring , kraftnät , transport och telekommunikationer .
jag vill framhålla att det interregionala samarbetet bidrar till att ansluta de lokala och regionala myndigheterna till den europeiska integrationsprocessen .
vi måste nämligen främja ett aktivare deltagande av de lokala och regionala myndigheterna när det gäller gemenskapsinitiativen , samtidigt som vi tar hänsyn till att de regionala och lokala myndigheterna ofta har mycket begränsad samarbetskapacitet på grund av mångfaldiga rättsliga ramar och utvecklingsnivåer på ena eller andra sidan av samma gräns .
inom ramen för det gränsöverskridande samarbetet bör vi lägga större vikt vid att förbättra driftsvillkoren för sysselsättningsskapande små och medelstora företag .
på samma sätt och mot bakgrund av att femtio procent av arbetslösheten är strukturell arbetslöshet bör de medel som ställs till förfogande från interreg vara tillräckligt stora för att komplettera nationella sysselsättningsfrämjande åtgärder .
mer konkret kan sägas att den gränsöverskridande rörligheten omöjliggörs , bromsas och blir problematisk på grund av hinder , som alltför ofta är anknutna till skattesystemet ( dubbelbeskattning ) och det sociala trygghetssystemet .
jag önskar att de projekt som ingår i programmen skall bidra till att finna lösningar på dessa problem och ge ett konkret innehåll åt den fria rörligheten för arbetstagare , en princip som i min region väger tungt !
interreg-anslagen bör också bidra till att inrätta ett europeiskt forskningsområde .
slutligen och framför allt finns det mycket stora förväntningar i regionerna på detta initiativ , eftersom kommunerna som inte är stödberättigade till mål 2 hoppas bli kompenserade tack vare interreg !
det är således viktiga saker som står på spel : införlivandet av gränsområdena kommer att utgöra en väsentlig faktor när den framtida europeiska regionalplaneringspolitiken utarbetas !
jag hoppas att var och en är lika medveten om det som f. decourrière som jag gratulerar !
. ( fr ) gemenskapsinitiativet interreg är en olycksdiger beståndsdel i den europeiska regionalpolitiken .
denna politik som till ytan verkar generös eftersom den officiellt är avsedd för att hjälpa områden i svårigheter är en narrarnas marknad för de franska skattebetalarna .
frankrike som bidrar med 17 procent av den europeiska budgeten , får bara 8 procent av de regionala strukturfonderna .
mellan 1994 och 1999 fick våra regioner genomsnittligen 15,4 miljarder franc per år , men de kommer bara att få 14,7 miljarder mellan åren 2000 och 2006 .
min region , nord-pas-de-calais , kommer att särskilt beröras , eftersom franska hainaut förlorar mål 1-stöden .
en oberättigad indragning i ett område vars främsta verksamheter har förstörts genom frihandelspolitiken i europa .
den europeiska regionalpolitiken stärker också bryssels centralregering , med vilken de regionala myndigheterna uppmanas förhandla direkt om användningen av strukturfonderna .
det är regionernas europa , regioner som inte har samma kraft som våra nationer och lätt kommer att foga sig efter bryssel .
interreg-initiativet som tillkom 1990 för att förbereda - jag citerar : &quot; gränsområdena till ett europa utan gränser , således utan nationer , passar mycket väl in i denna filosofi &quot; .
decourrière framför emellertid kloka reflexioner då han pekar på brysselteknokraternas brister .
dessa kommer i synnerhet att leda till ett försenat genomförande av interreg iii och således finansiella förluster för mottagarområdena .
vi är också ense med honom om att begära mer uppmärksamhet åt små och medelstora företag och naturligtvis vägra ta hjälp av ett externt tjänsteföretag .
det är sådana metoder som ligger bakom den föregående kommissionens korruptionsaffärer .
dessa punkter , som innehåller sunt förnuft och som vi har röstat för , rättar dock inte till den eurofederalistiska filosofi som präglar gemenskapsinitiativen , i synnerhet interreg .
därför röstade nationella fronten emot betänkandet .
. ( fr ) europaparlamentet har gett sin åsikt om kommissionens riktlinjer rörande gemenskapsinitiativet interreg om gränsöverskridande , transnationellt och interregionalt samarbete .
jag vill försvara ett ändringsförslag som ingavs av min grupp om frågan om detta initiativs havsdimension .
det handlar inte om att åter oroa sig för atlantbågens framtid utan om nödvändigheten att införliva principen om havsgränser i avdelning a rörande det gränsöverskridande samarbetet .
i europeiska kommissionens riktlinjer finns det inte många havsområden som är stödberättigade till interreg iii a. ändringsförslagen till betänkandet decourrière går mot en &quot; havsinriktning &quot; av interreg .
denna utveckling är viktig och bör fortsätta eftersom det är unionens framtid som står på spel .
jag känner till europeiska kommissionens motstånd i frågan . den framförde det vid samtalet i november om framläggandet av interreg iii .
men jag vill påpeka följande : att förhindra ett erkännande av havsgränserna betyder att man förnekar att det finns ett område som är potentiellt rikt på projekt och innovationer .
ett enda exempel : det så kallade &quot; keltiska &quot; området som omfattar områdena bretagne i frankrike , cornwall och devon i förenade kungariket , cork och waterfold i irland är ett område som har en närekonomi grundad på beroende av fiskerisektorn och betydelsen av lantbruket samt privilegierade kulturella och vänskapliga band ( vänorter ) .
interreg iii , avdelning a , skulle göra det möjligt för dessa områden att föra fram ett antal strukturprojekt som är nödvändiga för utvecklingen av små och medelstora företag samt för teknisk forskning och utveckling genom kunskapsöverföring .
det skulle således vara önskvärt att europeiska kommissionen kan delta i genomförandet av infrastrukturer för hamnar och flygplatser för förbindelserna mellan regionerna .
denna politik skulle således få stora ekonomiska konsekvenser för fisket i bretagne eftersom fisken skulle kunna landsättas på framskjutna irländska baser för att därefter skickas hem till livsmedelsföretagen i bretagne .
införandet av havsgränsen i avdelning a skulle göra det möjligt att äntligen erkänna ett enda ekonomiskt och stort område i västra randområdet inför europeiska unionens kontinentala förskjutning .
det skulle vara att visa respekt för dessa yttersta randområden som oroar sig en aning inför utvidgningen mot öster .
havsvärlden har en stor potential .
vi får inte åsidosätta den i gemenskapens nydanande pilotprogram som gör det möjligt att fastställa europas nya geografiska och ekonomiska karta .
( da ) det europeiska projektet startade som ett samarbete mellan stater .
detta samarbete har säkrat freden och stabiliteten i vår del av europa i över 50 år .
som ett resultat av de ekonomiska och politiska framgångarna i vår del av världen , som bl.a. eu är ett bevis på , och i och med den allt större spridningen av våra västliga värderingar , har konkurrensen på världsmarknaden vuxit kraftigt under de senaste årtiondena .
denna konkurrens skall eu vara redo att möta .
det kan vi bara göra genom att intensifiera samarbetet inom gemenskapen .
här handlar det inte om en större integration av länderna i form av en federation , utan om att utnyttja våra ekonomiska möjligheter över gränserna .
projekt som gör det möjligt att bygga ekonomiska tillväxtcentrum på gemenskapsnivå , som kommer att kunna anta utmaningen från våra konkurrenter på det globala planet .
jag välkomnar därför en fortsättning på programmet .
( fr ) betänkandet av decourrière saknar inte goda egenskaper ; denna lika tydliga som uttömmande presentation av interreg-initiativet och dess roll för att bryta gränsregionernas isolering ställer sig , i punkt 16 , på de små och medelstora företagens sida .
med min kollega dominique souchet , som är insatt i denna fråga , har jag ingivit fem ändringsförslag som framhåller de små och medelstora företagens och hantverkarnas roll inom ramen för interreg , betydelsen av samarbete mellan företag och kravet på att ekonomiska och sociala partner skall vara delaktiga i utformningen och genomförandet av programmen . dessa ändringsförslag har antagits enhälligt , vilket gläder mig .
men den franska delegationen i vår grupp kan inte acceptera att kommissionen och den federalistiska klanen avleder interreg-initiativet från dess syfte , för att ytterligare försvaga nationernas politiska roll .
vi avser inte att låta bryssel ta hand om medlemsstaternas regionala fysiska planering , vilket skäl l i betänkandet antyder .
vi begär bara en sak från kommissionen : att den nöjer sig med att se till att genomförandet av gemenskapens politik inte hotar en balanserad fysisk planering .
den gemensamma jordbrukspolitiken och emu : s skadliga effekter för balansen mellan olika regioner och framför allt för vitaliteten i de mest avlägsna och glesbefolkade landsbygdsregionerna , visar att en sådan ambition är allt annat än ett latmansgöra .
därför kan vi inte godkänna utvecklingen av området iiic i gemenskapens initiativ , ett område som genom att uppmuntra samarbetet mellan regionerna under kommissionens ansvar håller medlemsstaterna vid sidan om .
den förtjusning som uttrycks för område iiic blir desto märkligare då föredraganden i sin motivering själv erkänner att &quot; utkastet till riktlinjer &#91; innehåller &#93; inga uppgifter om eventuella samarbetsområden &quot; ( s.16 ) och att &quot; ansvaret är &#91; ... &#93; oklart &quot; ( p.17 ) .
att under sådana omständigheter kräva ytterligare medel för detta avsnitt , som i punkt 20 , är ännu ett av de lika oansvariga som ideologiska överbud som kammaren är sin vana trogen .
låt oss till sist konstatera det felaktiga i den vilja som uttrycks såväl i kommissionens dokument som i betänkandet av decourrière : att interreg skulle användas för freden och återuppbyggnaden på balkan . jag tror inte att strukturfonderna skall utnyttjas för att reparera de skador som amerikanerna har åsamkat serbien i samband med de både brottsliga och ineffektiva bombningarna .
det är washingtons sak och inte vår , att ta på sig ansvaret för en konflikt som de utlöste för att tjäna sina egna intressen .
därför har den franska delegationen i vår grupp inte kunnat stödja decourrièrebetänkandet . vi har valt att avstå vid den slutliga omröstningen .
betänkande ( a5-0025 / 2000 ) av procacci
herr talman ! jag röstade för procaccis betänkande om landsbygdsutveckling , inte bara för att jag instämmer i huvuddragen i leader-programmet utan också för att det är den andra sidan av urban-programmet , som vi talade om tidigare .
precis som de äldre i städerna är mycket ensamma börjar de äldre på landsbygden bli den enda kvarvarande befolkningen , eftersom de unga flyttar till städerna : de dras till ljusen , till barerna också , och landsbygden töms .
jag tror alltså att det är mycket viktigt att detta projekt inom europeiska unionen får stöd av alla och byggs ut ytterligare .
. ( pt ) det gemensamma initiativet leader + , även om det är en fortsättning på tidigare initiativ , uppvisar en del besynnerligheter .
först och främst halveringen av de tillgängliga anslagen , trots att perioden förlängts .
likväl inkluderas nya mål , till exempel finansieringen av natura nätverk 2000 , och landsbygden blir ett annat valbart alternativ .
trots att det här gemenskapsinitiativet avser landsbygdens tillväxt tar man inte samstämmigt upp jordbruket och jordbruksproduktionen , och detta är inte rimligt .
ingen landsbygd utan jordbruk , vilket gör att vilken strategi som helst för landsbygdens tillväxt måste baseras på jordbrukets endogena potential , oaktat andra aktiviteters större eller mindre tillväxt för att hindra landsbygdens desertering .
därför menade vi att det var så viktigt att förbättra betänkandet med de förslag som vi lade fram om att jordbruksaktiviteterna och lantbrukarna uttryckligen borde inkluderas i strategin för landsbygdens tillväxt , och att man borde ansöka om större anslag så att man kan fortsätt med programmet på de orter som tidigare inkluderats samt ta det nya programmet , som skall fortsätta att privilegiera de minst gynnade områdena , i försvar .
min inställning till leader hänger samman med min inställning till eu : s jordbrukspolitik över huvud taget .
såväl leader i som leader ii , vilka genomförts under 1990-talet , har ingått i den nya gemensamma jordbrukspolitik som tillämpats allt sedan revideringen 1992 och har tillsammans med andra åtgärder utgjort den s.k. andra pelaren i eu : s politik för landsbygdsutveckling .
deras verkliga syfte har varit att förringa och skyla över de katastrofala följderna av den nya gemensamma jordbrukspolitiken och att vilseleda de små och medelstora jordbruken , och de har inte haft till syfte att utveckla landsbygden och att behålla jordbruksbefolkningen på landsbygden , vilket man så hycklande brukar påstå .
detta framgår av det faktum att jordbruksinkomsterna och sysselsättningen har minskat mycket hastigt i de områden där dessa initiativ har tillämpats , vilket lett till allt snabbare avfolkning av dessa områden . grekland är ett betecknande exempel .
som mål 1-land omfattades grekland i sin helhet av gemenskapsinitiativen från leader . samtidigt minskade sysselsättningen inom jordbruket med 2,3 procent under perioden 1994-1999 , medan jordbruksinkomsterna minskade med 15,2 procent .
jag anser att leader + kommer att vara effektivare än leader i och ii av följande orsaker .
de verkliga målen för leader + är de samma som för leader i och ii . dvs. att mildra och skyla över de negativa effekterna av den gemensamma jordbrukspolitik som kommer att tillämpas inom ramen för agenda 2000 .
men denna gemensamma jordbrukspolitik är sämre än den föregående och dessutom har den ett sämre utgångsläge , eftersom revisionen av den gemensamma jordbrukspolitiken 1992 och gatt-avtalet 1995 har lett till betydande problem och svårigheter för jordbruksekonomin .
urvalskriterierna och de verksamheter som finansieras genom leader kan i bästa fall lindra enstaka mindre viktiga landsbygdsproblem , men i värsta fall urartar de till offentliga utgifter som bara tjänar till att döva samvetet .
programmen leder inte till någon allsidig utveckling av de utvalda områdena och de leder inte heller till nya , stadigvarande arbeten på landsbygden , för de flesta verksamheterna har inte någon produktiv inriktning .
de verkliga anslagen till leader + är mindre än anslagen till leader ii , trots en ökning med 15 procent ( från 1775 miljoner euro för leader ii till 2020 miljoner euro för leader + ) .
och detta beror på att ökningen med 15 procent är nominell och inte reell , eftersom den genomsnittliga årliga inflationen inom gemenskapen under dessa år uppgår till ungefär 2 procent .
leader + pågår ett år längre än leader ii .
till leader + kan man föra alla eu : s regioner , medan leader ii omfattade mål 1-regionerna och vissa regioner inom mål 5b och 6 .
men jag vill påpeka att även om de reella anslagen till leader + var högre , så skulle gemenskapsinitiativet ändå vara ineffektivt , eftersom den jordbrukarfientliga inriktningen av den gemensamma jordbrukspolitiken inom ramen för &quot; agenda 2000 &quot; inte kan vare sig kompenseras eller mildras av sådana program som i många områden endast syftar till att skyla över , att vilseleda och att döva samvetet .
jag motsätter mig många av åsikterna i betänkandet .
jag vill ännu en gång påpeka de negativa förändringarna i den gemensamma jordbrukspolitiken ( 1992 - agenda 2000 ) .
jag anser att leader + inte kommer att bidra till en verklig lösning av landsbygdens problem , med allt svårare förhållanden för jordbruket , som ju har varit och bör vara den viktigaste samhällsekonomiska näringsgrenen på landsbygden .
jag kommer för min del att informera jordbrukarna om syftet med dessa program .
jag kommer att verka för att de skall utnyttjas på bästa tänkbara sätt utan att slösas bort och , framför allt , kommer jag att verka för att utveckla jordbrukarnas kamp mot den katastrofala gemensamma jordbrukspolitiken , som utarmar dem och leder dem till ekonomisk bankrutt , samtidigt som landsbygden avfolkas .
om man inte avskaffar denna gemensamma jordbrukspolitik , finns det nämligen inget program som kan garantera att de små och medelstora jordbruken överlever och att landsbygden vitaliseras socialt och ekonomiskt .
. ( fr ) samtliga ledamöter i gruppen unionen för nationernas europa har röstat för nästan allt i betänkandet av vår kollega procacci rörande gemenskapsinitiativet leader + .
vi har emellertid ändrat det förslag till betänkande som hade godkänts av utskottet för jordbruk för att klarlägga vissa punkter varvid gemenskapsinitiativet kunde göras mer operativt .
det verkar för oss väsentligt att i synnerhet förenkla de administrativa och finansiella förfaranden som visade sig bli för tunga och långsamma inom ramen för initiativet leader ii .
det verkar också nödvändigt att säkra att bättre hänsyn tas till de lokala aktörernas utvecklingsprioriteringar och att inte utdelningen av fonderna leader + bara begränsas till jordbruksområden med låg befolkningstäthet .
i ändringsförslag 10 , som jag har ingett på min grupps vägnar , hänvisas till begreppet &quot; ekonomisk och social sammanhållning &quot; i stället för &quot; regionalplanering &quot; eftersom europeiska unionen inte har erkänd befogenhet på området .
i ändringsförslag 11 ersätts termerna &quot; statlig eller kommunal administration &quot; med &quot; samtliga offentliga förvaltningar &quot; .
de lokala åtgärdsgrupperna bör visserligen utgöra en balanserad enhet som är representativ för partner från olika socioekonomiska miljöer i området men på beslutandeplanet bör i själva verket samtliga offentliga förvaltningar ( kommuner , län , regioner och stater ) företrädas i sin helhet vilket nivå de än har .
föredragandens formulering var således alltför inskränkande , enligt vår åsikt .
vad beträffar ändringsförslag 12 uppfyller det förväntningarna i europaparlamentets utskott för regionalpolitik .
det inbegriper den nödvändiga samordningen mellan leader + och gemenskapsprogrammen för samarbete och partnerskap , såsom interreg , phare , sapard eller meda .
på europeiska unionens , kandidatländernas och efta : s medlemsstaters territorium kan det finnas interna förbindelser mellan de olika gemenskapsinitiativen .
man måste komma ihåg att de verkliga prioriteringarna för den europeiska världsdelen är att införa en operativ nivå inom europeisk ram och inte inom en global ram , såsom föredraganden föreslår .
skapandet av organisationer liknande lokal åtgärdsgrupper ( gal ) kan med fördel uppmuntras av europeiska unionen , naturligtvis förutsatt att motsvarande kostnader bestrids av de olika parterna .
vi ställer oss i grund och botten naturligtvis positiva till gemenskapsinitiativet leader + .
vi måste komma ihåg att vid konferensen om landsbygdsutveckling som hölls i cork den 7-9 november 1996 definierades landsbygdsutveckling såsom en av europeiska unionens prioriteringar eftersom det är av största vikt att bevara vårt jordbruks och hela landsbygdsstrukturens ( infrastrukturer , offentliga och privata tjänster ... ) integritet .
i det sammanhanget har vi i utskottet beklagat avsaknaden av anslag för landsbygdsutveckling och stött de ändringsförslag som begär en ökning av budgeten för detta gemenskapsinitiativ , så att det kommer i jämvikt med de tidigare initiativen leader i och leader ii .
jämfört med det senare initiativet som hade begränsad giltighetstid på sex år , är den anslagna budgeten för leader + femtio procent lägre för en period av sju år .
det är inte godtagbart med tanke på den betydande landsbygdsutvecklingen och konsekvenserna för jordbrukarna av pris- och stödsänkningarna enligt den planerade reformen av den gemensamma jordbrukspolitiken till följd av berlinavtalen .
bland de prioriterade kriterier som kommer att införas på europeisk nivå för att möjliggöra lokala anmälningar bör slutligen särskild uppmärksamhet ägnas åt de projekts kvalitet och originalitet som redan uppburits av gal inom ramen för initiativet leader ii men som inte kunnat slutföras på grund av tidplanen och de omständliga planerade förvaltningsåtgärderna .
nästa punkt på föredragningslistan är betänkande ( a5-0015 / 2000 ) av graefe zu baringdorf för utskottet för jordbruk och landsbygdsutveckling om förslaget till rådets direktiv om ändring av direktiv 70 / 524 / eeg om fodertillsatser ( kom ( 1999 ) 388 - c5-0134 / 1999 - 1999 / 0168 ( cns ) ) .
herr talman , herr kommissionär ! har regleringen av fodertillsatser att göra med konkurrens eller med konsumentpolitik ?
för kommissionen och utskottet för rättsliga frågor är det en fråga om konkurrens .
säkerligen måste vi ta hänsyn till djurfoderindustrins konkurrenskraft när föreskrifterna för ämnen som tillåtits före och efter 1988 harmoniseras .
det bör förhindras att priset på djurfoder höjs , och därför bör doyles ändringsförslag 4 och 5 stödjas .
men i första hand är det , som graefe zu baringdorf formulerat det i sitt betänkande , en konsumentpolitisk fråga .
livsmedelssäkerheten måste ha absolut prioritet i alla diskussioner om djurfoder .
när vi talar om öppenheten i näringskedjan , så gäller det från dynggrepen till bordsgaffeln , och därför börjar alltså konsumentskyddet med djurfodret .
antibiotika , tillväxtbefrämjande medel och genetiskt modifierade organismer hamnar ändå till slut i människans näringskedja .
som en konsekvens av dioxinskandalen blev det klart för oss alla att vi äntligen måste ta oss ur detta mörka hörn . regleringen av fodertillsatserna är ett steg i rätt riktning .
enligt artikel 152 i eg-fördraget är vi ålagda att undanröja sådana orsaker som kan hota människans hälsa . betoningen ligger entydigt på orsaker .
helt konsekvent måste vi stänga av de ursprungliga källorna till skadliga ämnen - nämligen skadliga fodertillsatser .
i annat fall , anser jag , laborerar vi med symptomen , men vi bekämpar inte orsakerna .
befolkningen är mycket kritisk i synnerhet när det gäller användning av gmo .
vi måste ta hänsyn till befolkningens ökande känslighet beträffande gmo , och reglera användningen i djurfoder i enlighet med detta .
för det första : om en tillsats består av genetiskt modifierade organismer , eller om den innehåller sådana organismer , får denna tillsats bara tillåtas om den är ofarlig för människans hälsa och för miljön .
för det andra : det är förnuftigt att analogt med bestämmelserna i lagen om avyttring av utsäde , vilket även föredraganden har berört , utfärda föreskrifter för genetiskt modifierade fodertillsatser .
och för det tredje : för att få en öppen konsumentpolitik behöver vi en märkning av genetiskt modifierat djurfoder .
denna entydiga innehållsdeklaration för djurfoder möjliggör alltså en dubbel beslutandefrihet , både för den som använder djurfoder och för den senare konsumenten .
beslutet bör ligga hos den myndigförklarade medborgaren , anser jag .
vi talar alla om de skandalöst pungslagna medborgarna , som har förlorat förtroendet för livsmedelssäkerheten .
med en konsekvent reglering av fodertillsatserna kan vi nu bidra väsentligt till att återvinna förtroendet .
därför är jag alltså mycket spänd på att få höra ert svaromål vad gäller våra ändringsförslag .
alltså kommer vi naturligtvis att rösta så att vi eventuellt skickar tillbaka förslaget till utskottet .
herr talman , kära kolleger ! föreliggande förslag till ändring av direktivet om fodertillsatser från år 1970 är det första i en hel rad förslag när det gäller djurfoder .
vi kommer alltså under de närmaste månaderna här i parlamentet att diskutera ytterligare några .
att denna fråga har central betydelse bevisar den stora uppmärksamhet som den europeiska allmänheten har skänkt skandalerna med dioxin , antibiotika , slam från reningsverk osv. det handlar här alltså om en viktig beståndsdel i skyddet av allmänhetens hälsa .
därför anser vi att artikel 152 skall användas som rättslig grund och inte artikel 37 , som kommissionen har föreslagit .
den ändring som kommissionen har föreslagit , nämligen lika behandling av de tillsatser som godkänts efter respektive före den 31 december 1987 , är oomtvistad , och har vårt fulla stöd .
utskottet för jordbruk och landsbygdens utveckling har dock enhälligt gjort några viktiga ändringar i kommissionens förslag .
de av kommissionen föreslagna bestämmelserna medför risk för monopolbildning vid saluförandet av vissa tillsatser .
förslagsrätt medges endast dem som erhållit det ursprungliga godkännandet , men utesluter de företag som senare har fått ett godkännande .
en sådan monopolbildning , som exempelvis skulle kunna leda till en höjning av priset på djurfoder , bör vi förhindra genom att ge ett preliminärt godkännande till alla företag som den 1 april 1998 saluförde ett visst ämne .
detta skall sedan gälla tills den förnyade utvärderingen har avslutats .
den viktigaste ändringen gentemot kommissionens förslag gäller dock det av föredraganden rekommenderade inkluderandet av bestämmelser om genetiskt modifierade organismer i direktivet om tillsatserna . han har här utgått från den kompromiss som parlamentet och kommissionen kommit överens om beträffande godkännande av genetiskt modifierade organismer utanför utsättningsdirektivet .
denna utgör redan grundvalen för godkännandet av genetiskt modifierade organismer .
därför är det bara logiskt och i enlighet med de bestämmelser som vi redan har godkänt på andra områden - jag kan bara nämna skogsodlingsmaterial - att även i föreliggande fall föreskriva bestämmelser om genetiskt modifierade fodertillsatser .
här spelar i synnerhet märkningen av genetiskt modifierade tillsatser en viktig roll .
å ena sidan medger den att jordbrukaren kan fatta ett medvetet beslut om huruvida han vill använda sådant djurfoder eller inte , och å andra sidan blir det möjligt för konsumenten att avvisa livsmedel som framställts på basis av genetiskt modifierade organismer .
avslutningsvis också ett hjärtligt tack från vår grupp till föredraganden , som lagt ner mycket arbete på detta .
jag tror vi kan vara nyfikna på att få höra vad byrne kommer att säga .
detta betänkande handlar mer om formerna , dvs. hur tillsatsämnen skall godkännas , och något mindre om vilka de är och hur de fungerar .
jag måste få ta tillfället i akt att understryka hur viktigt det är att alla dessa direktiv i fortsättningen behandlas enligt förfarandet i artikel 152 , eftersom både livsmedelssäkerhet och miljöfrågor kräver en sammanhållen politik , en helhetssyn .
vi kan inte göra som vi gjort hittills , dvs. ta varje detalj för sig och ofta först när skadan redan är skedd .
föredraganden har betonat prövning och märkning av gmo i fodertillsatsen .
jag skulle än en gång vilja tala om antibiotika .
förvisso är fem av de nio antibiotika som ursprungligen var tillåtna i foder i dag förbjudna , men det är oerhört viktigt att vi förbjuder även de sista fyra , inte bara för folkhälsans , utan även för djurens skull .
vi har kommit så långt att vi känner till antibiotikaresistensens oerhörda hot mot folkhälsan , framför allt för småbarn .
i många medlemsstater kan man redan bevisa att missbruket i djurhållningen är helt onödigt .
det finns flera länder som för länge sedan har fasat ut foderantibiotika , och det finns några som är på väg att göra det med lyckat resultat .
försiktighetsprincipen , som vi talar mycket om , har vi för länge sedan gått förbi , när det handlar om antibiotika .
det finns emellertid ytterligare en princip i miljöarbetet som är viktig , nämligen utbytesprincipen .
jag skulle vilja säga något kort om coccidiostatika .
det är ett tekniskt antibiotikum , som inte är absolut nödvändigt .
det finns ersättningsmedel . det går att vaccinera kycklingar .
det kostar visserligen litet mer , men är ofarligt för miljön .
i dag åker coccidiostatika ut med gödseln på åkern .
därmed hamnar det i vattnet som ju faktiskt är vårt viktigaste livsmedel .
herr talman , herr kommissionär , mina kära kolleger ! betänkandet om fodertillsatser avser ett teknisk-ekonomiskt problem för att återställa konkurrensjämvikt mellan de olika fodertillsatserna och mellan tillsatsernas producenter .
men nu efter den allvarliga dioxinkrisen som drabbade belgien och andra europeiska länder förra sommaren kan man inte nöja sig med att diskutera om en enkel konkurrensfråga .
en gång i tiden , även om det gick mer obemärkt förbi allmänheten , upptäckte nämligen kommissionens vetenskapliga experter industriella kalkrester fulla med dioxin i pressade citrusfrukter som importerats från brasilien .
därför är det tid att redovisa samtliga beståndsdelar i den kedja som deltar i tillverkningen av foder för avkastningsdjur .
vi kan i förbigående konstatera , och det är en skandal , att problemet är mycket mindre allvarligt när det gäller foder för våra hundar , katter och övriga husdjur .
är det på grund av den vilda och globaliserade konkurrens som denna sektors industrier ägnar sig åt som den har omvandlats till en återvinningssektor för avfall från livsmedelssektorn ?
ett så allvarligt ämne kan inte begränsas till en teknisk debatt även om det ju är det direktiv som begränsar tillståndet för antibiotika och andra tillväxtfaktorer .
de försiktighetsåtgärder som vi gör oss beredda att vidta för djurfoder bör också tillämpas i fråga om foder till lantdjur , just de djur som vi återfinner på tallriken .
såsom det med kraft betonas i betänkandet är märkning en absolut nödvändighet så att varje jordbrukare i sitt företag känner till samtliga ingredienser som ingår i det foder som han avser att ge till sin besättning .
han bör också veta om genetiskt modifierade organismer , gmo , har trängt in i hans proteinkornspåse . dessa beståndsdelar kan potentiellt utgöra en folkhälsorisk .
genom försiktighetsprincipen har vi i varje fall fått krav om en tydligt angiven spårbarhet på alla nivåer vid saluföringen av dessa produkter .
men före märkningen måste tydliga regler införas .
man måste ställa enkla frågor såsom frågan om det verkliga syftet med användning av djurfoder .
om vi betraktar alla problem som det har åsamkat oss ur etisk synpunkt och sanitär synpunkt , måste vi nu ställa oss frågan om själva användningen .
det kapitel i vitboken om livsmedelssäkerhet , som behandlar djurfoder , bör i det avseendet tjäna som grund för arbetet med att gå långt bortom de enkla saluföringsfrågorna .
kommissionen har vid flera tillfällen använt följande exempel : &quot; från grepen till gaffeln &quot; . vår kollega i ppe betonade det nyss .
det är en god formulering , men vi måste också ge den mening . och för att ge den mening måste vi behandla såväl problemen med djuren som problemen med konsumenternas hälsa .
därför är det viktigt att godkänna ändringsförslag 2 till skäl 4 , som gör det möjligt att undvika risk för monopol , om de bolag som först fick tillstånd att saluföra en tillsats skulle förbli de enda som kunde utnyttja det under omvärderingsperioden .
men ändringsförslag 4 och 5 till den nya artikel 2 a måste framför allt godkännas , eftersom de gör det möjligt att tydligt utpeka tillsatser som är genetiskt modifierade för att användarna skall kunna fatta beslut med full sakkännedom .
herr talman , mina damer och herrar ledamöter ! användningen av tekniskt avancerade tillsatser inom djurfoderbranschen kräver detaljerad information från aktörerna - och det är som bekant ganska många - om deras insatser , för att man skall förhindra metoder som bryter mot gemenskapsrätten .
det befintliga direktivet om fodertillsatser kan inte ensamt åstadkomma detta .
det kommer att följas av andra direktiv , och jag anser att de är på rätt plats i utskottet för jordbruk och landsbygdens utveckling .
innan kött , mjölk , bröd och andra produkter försäljs över disk kommer djurfoder och tillsatser att struktureras , blandas , mixas , skäras sönder och transporteras upprepade gånger .
kampen bland djurfoderproducenterna för att uppnå största marknadsandel innebär , på samma sätt som inom livsmedelsproduktionen , många problem .
de negativa följderna känner vi till , de positiva vet vi mindre om .
jag är fast övertygad om att hälsan för de europeiska konsumenterna i den ekologiska kedjan bäst kan skyddas genom att livsmedel och djurfoder produceras inom regionen och för regionen .
men detta kräver ytterligare arbete .
herr talman ! får jag börja med att gratulera föredraganden , graefe zu baringdorf , för hans betänkande .
det avspeglar åsikterna och oron hos alla eu-medborgare över frågor som rör livsmedelssäkerhet och livsmedelskvalitet .
tidigare händelser under ett antal år har förvisso skapat en medvetenhet och farhågor om det verkliga hotet mot livsmedelssäkerhet och folkhälsa .
den snabba insats som görs av detta parlament måste av alla medborgare anses som deras största garanti för framtiden för ni har lagt fast en dagordning om livsmedelskvalitet som medlemsstaterna måste rätta sig efter .
men även på detta viktiga förvaltningsområde visar parlamentet sitt åtagande om subsidiaritet genom att uppmuntra medlemsstaterna att ta på sig sitt ansvar .
i agenda 2000 har vi enligt min åsikt prioriterat politikområden som direkt berör medborgarna : livsmedelssäkerhet , vattenkvalitet , miljöskydd och utveckling av landsbygden .
om vi fullföljer denna dagordning med engagemang och hårt arbete kommer de första åren av det nya millenniet att bli en milstolpe för genomförandet av en politik som är inriktad på människorna och som väldigt mycket speglar gemenskapens behov .
jag välkomnar i synnerhet de föreslagna nya och strikta tillståndsförfarandena för tillsatser i djurfoder .
de som upptäcks bryta mot dessa måste behandlas strängt .
jag gratulerar den nye kommissionären , byrne , som ansvarar för livsmedelssäkerhet .
han har en tung uppgift men har agerat snabbt och effektivt på kraven från denna kammare , liksom på konsumenternas oro .
jag är särskilt glad att mitt eget land , irland , ligger i frontlinjen med genomförandet av nya livsmedelsföreskrifter grundade på principen om spårbarhet .
detta kommer att göra ön irland till ett framstående centrum i framtiden när det gäller livsmedelsproduktion .
jag skulle också vilka gratulera föredraganden som har gjort ett utmärkt arbete och framför allt glädja mig åt den enhällighet som har rått på gruppnivå om detta ärende .
det är således planerat att kommissionen skall byta ut de befintliga tillstånden mot tillstånd knutna till de ansvariga för saluföringen av tillsatserna genom en förordning och att dessa byten skall göras på samma gång i fråga om alla berörda tillsatser .
vi måste återställa en sammanhållen rättslig ram .
kommissionen föreslog att införa en rättslig grund från och med oktober 1999 i direktiv 70 / 524 / eeg för att ersätta tillstånden .
vi måste emellertid se till att inte skapa snedvridningar av konkurrensen såsom kindermann och auroi påminde om .
jag tror att vi också tydligt måste identifiera de genetiskt modifierade tillsatserna i djurfoder för att göra det möjligt för och garantera för slutkonsumenten att han kan välja gmo-fri mat eller mat baserad på gmo .
konsumenten bör få behålla sin beslutsfrihet med full sakkännedom .
detta förslag har ingen finansiell inverkan på gemenskapens budget , herr kommissionär .
därför behöver vi för livsmedelssäkerheten en total öppenhet för producenterna och konsumenterna .
jag är övertygad om att kommissionen kommer att kunna följa föredraganden som , vill vi påminna om , har uppnått enhällighet i utskottet för jordbruk och landsbygdsutveckling .
herr talman ! sedan bse först dök upp har vi här i kammaren alltid sagt att djurfodret är en av de första och viktigaste beståndsdelarna för en säker produktion av livsmedel , för att skydda konsumenternas hälsa .
därför gläder det oss att kommissionen lägger fram ett förslag om fodertillsatser .
utskottet , som jag här talar för , nämligen utskottet för miljö , folkhälsa och konsumentskydd , beslutade i december - förutsatt att ordföranden i utskottet för jordbruk och landsbygdens utveckling i egenskap av föredragande skulle utarbeta ett sådant bra betänkande - att vi kan avstå från ett yttrande .
trots detta vill jag säga ett par saker och ta ställning till några punkter .
först kanske något om den rättsliga grunden .
även om vi i parlamentet har en ny arbetsordning - och det mycket väl kan hända att det med den mycket ambitiöse ordföranden i utskottet för jordbruk allt oftare kan uppstå tvister mellan utskottet för jordbruk och utskottet för miljö när det gäller ansvarsområdet för lagstiftningen - är trots detta en sak helt klar för mig när det gäller sådana konflikter : sammanhållningen i parlamentet är avgörande , och den rättsliga grunden i en fråga är avgörande för mig .
därför - det måste jag säga er , herr byrne - fördömer jag den rättsliga grund som valts .
om den endast är en traditionell rättslig grund som övertagits från de tidigare direktiven , då är det fel att bibehålla den .
amsterdamfördraget säger helt klart : när det gäller människors hälsa skall artikel 152 väljas som rättslig grund , och jag måste här säga till utskottet för rättsliga frågor och den inre marknaden i vår egen kammare : det räcker helt enkelt inte att titta på kommissionens förslag och säga att det inte står någonting i det om hälsa och konsumentskydd , alltså handlar det inte heller om hälsa och konsumentskydd .
därför kommer min grupp - som kindermann redan sagt - i morgon att rösta för en ändring av den rättsliga grunden , och jag hoppas att de andra grupperna i kammaren också kommer att göra det .
herr byrne , jag ber er för öppenhetens och det goda samarbetets skull att anta och rösta för en ändring av den rättsliga grunden .
om vi nämligen inte gör det , utan hörsammar utskottet för rättsliga frågor , skulle vi öppna dörren för manipulation .
då tillåter vi nämligen kommissionen att välja den rättsliga grunden , så att politiken för folkhälsan helt enkelt inte nämns i texten , och då är det plötsligt fråga om artikel 37 .
låt mig helt kort också säga något om de två andra punkterna : beträffande genetiskt modifierade organismer i djurfoder får det inte vara så att man hänvisar till vertikal lagstiftning och säger att vi så småningom behöver en annan lagstiftning .
men den har vi för närvarande inte !
och så länge som vi inte har det , måste vi alltid när vi beslutar om lagstiftning också behandla genetiskt modifierade organismer , nämna dem särskilt och insistera på en märkning .
det har föredraganden gjort , och det är ett bra tips .
jag vill än en gång säga det som jag redan sagt många gånger : ja , jag vill att kommissionen gör upp förslag till en positivlista . vi kommer säkert sedan att diskutera och behandla den kontroversiellt i denna kammare , men vi behöver åtminstone ha ett förslag till en positivlista för fodertillsatser .
det är lika viktigt att vi har stränga hygieniska krav på produktionen av tillsatser och att det kontrolleras ordentligt i medlemsstaterna .
på båda områdena finns det fortfarande brister , och där har vi fortfarande mycket att göra .
herr talman ! jag vill gratulera föredraganden till hans betänkande .
detta är en fråga som vi utan tvivel skall överväga på nytt vid flera tillfällen i framtiden .
det som har hänt under de senaste åren har gjort oss uppmärksamma på de ofantliga problem som inte bara producenter av livsmedel utan även konsumenter kan vänta sig .
vi måste hitta en balans mellan dem .
vi måste lösa denna fråga eftersom det är viktigt att konsumenter återfår förtroendet för den mat de äter .
ett sätt att uppnå detta är att införa total insyn när det gäller märkningen .
genetiskt modifierade organismer ( gmo ) är den nya utmaningen för oss .
detta är något som människor är mycket oroade över och helt med rätta och jag själv delar denna oro .
men jag anser att vi inte skall tillåta vår oro över gmo överskugga vår oro över växtfrämjande ämnen i djurfoder eller antibiotika i foderblandningar .
i själva verket bör vi inte låta gmo skymma det faktum att kött- och benmjöl fortfarande ingår i djurfoder i många länder i europa .
en faktor bakom denna utveckling som har nämnts i denna debatt är konkurrensen - konkurrens mellan medlemsstater om kostnaderna för livsmedelsproduktionen .
detta är samtliga områden där vi måste säkerställa spelregler på samma nivå : livsmedel måste vara av samma standard i alla medlemsstater .
vi har haft dioxinskräckupplevelsen , bse och många andra problem .
huvudproblemet är av ekonomisk art , nämligen vem bär kostnaden ?
problemet är att kostnaden inte delas lika mellan konsumenten och producenten : producenten har tvingats bära alla kostnader .
vi behöver en rättvis fördelning av de extra kostnader som uppstår .
vi måste också se till att det livsmedel som importeras till europeiska unionen håller samma standard som inom europeiska unionen .
om vi inte bibehåller dessa standarder för importerade livsmedel kommer vi att möta större svårigheter i framtiden .
( en ) jag skulle först vilja tacka utskottet för jordbruk och landsbygdens utveckling och dess föredragande , utskottets ordförande , graefe zu baringdorf , för hans granskning av kommissionens förslag .
kommissionens förslag är som några av er sagt ganska teknisk .
ändå har den ganska enkla mål : att harmonisera förfarandena gällande tillstånd för fodertillsatser .
för närvarande skiljer sig handläggningen av tillstånd beroende på om ansökan lämnades före eller efter den 1 januari 1988 .
syftet med kommissionens förslag är att harmonisera förfarandena för att kunna garantera att inga sådana skillnader finns .
det föreslagna ändringsförslagets räckvidd är därför mycket begränsad .
fem ändringsförslag har lagts fram av parlamentet .
jag beklagar att kommissionen inte har möjlighet att godkänna dessa ändringsförslag trots det faktum att jag är helt medveten om uppfattningar och åtaganden hos parlamentet , utskottet för jordbruk och i synnerhet föredragande , graefe zu baringdorf , i dessa frågor .
jag skall ta upp vart och ett av de enskilda ändringsförslagen separat .
i det första ändringsförslaget föreslås en ändring av den rättsliga grunden för förslaget och att ersätta artikel 37 med artikel 152 .
jag vill endast påpeka att kommissionens förslag inte innehåller hänvisningar till hälso- eller konsumentskydd .
den föreslagna ändringen är teknisk och kan inte tolkas ha som primärt syfte att skydda folkhälsan .
jag konstaterar att parlamentets utskott för rättsliga frågor och den inre marknaden också godkänner att artikel 37 är den lämpliga rättsliga grunden .
jag vill påminna parlamentet om att i artikel 152 är hälsoskyddet det primära målet .
jag rekommenderar er de argument som anges i skrivelsen från utskottet för rättsliga frågor i vilken ståndpunkten fastslås med enligt min åsikt precision , tydlighet och med lovvärd kortfattad text .
ändringsförslag 2 och 3 syftar mycket längre än kommissionens förslag eftersom syftet med dem är att införa ytterligare bestämmelser om genetiskt modifierade tillsatser .
jag är den förste att gå med på att gmo är en mycket viktig fråga .
jag godtar och erkänner också att ett antal initiativ för att aktualisera eu-lagstiftningen på området gmo krävs .
detta tekniska ändringsförslag är emellertid inte det rätta instrumentet för att införa sådana initiativ .
kommissionen anser att det är för tidigt att ändra de nuvarande fastslagna bestämmelserna i direktiv 70 / 524 om genetiskt modifierade tillsatser i detta skede .
i stället är det lämpligt att vänta på utvecklingen i förbindelse med den gemensamma ståndpunkten om ändringsförslag till direktiv 90 / 220 , vilken just nu är under den andra behandlingen i parlamentet .
kommissionen planerar att gå mycket längre än vad som för närvarande föreslås av parlamentet i dess ändringar .
jag kan även försäkra parlamentet att jag skall se till att de relevanta bestämmelserna i direktiv 90 / 220 innefattas i förslaget om en omarbetning av direktiv 70 / 524 som kommissionen föreslog i vitboken om livsmedelssäkerhet som skall läggas fram för parlamentet innan juli månad 2001 .
jag kan också försäkra parlamentet att alla yttranden här i dag kommer att beaktas till fullo .
ändringsförslag 4 och 5 kan inte heller godkännas för att de ger obefogat företräde till imitationsprodukter genom att bevilja tillstånd att omsättas till och med innan en ansökan om tillstånd har ingivits .
kommissionen vidhåller att sådana ansökningar först skall bedömas i fråga om säkerhet och verkan innan tillstånd ges .
jag kan bara be er igen att lägga på minnet den tekniska formen i kommissionens förslag och att avvakta det verkliga förslaget till ett nytt direktiv om fodertillsatser för att ta itu med större frågor .
jag vill endast ta upp några av de specifika frågor som togs upp under debatten .
för det första , avseende synpunkter från herr graefe zu baringdorf , vill jag försäkra honom att vi kommer att ändra förfarandet för tillstånd till gmo tillsatser i tillsatsdirektivet 70 / 524 och inte i det nya foderdirektivet .
detta är ett direktiv som mer specifikt behandlar råmaterial snarare än tillsatser .
den text som parlamentet använde härrör från det direktiv som antogs 1998 .
men den vertikala lagstiftningen i direktiv 90 / 220 om hur man bedömer miljörisker i samband med gmo har förändrats sedan dess och håller fortfarande på att förändras .
det behandlas av parlamentet i en andra behandling .
jag tror att vi bör vänta på det slutliga resultatet gällande direktiv 90 / 220 och i synnerhet , artikel 11 .
man tog även upp frågan om detta förslag kunde skapa en risk för att monopol inrättades .
kindermann och auroi anspelade på detta .
jag vill endast ta upp några punkter i den frågan .
för det första har detta ärende funnits i stöpsleven sedan 1993 , så det har faktiskt inte överrumplat några andra råvaruproducenter .
varje sådan sökande kan i själva verket fortfarande lämna in en ansökan gällande sin speciella produkt .
ja vill också understryka att kommissionen aldrig har godkänt någon ansökan om tillstånd att använda gmo i tillsatser .
roth-behrendt berörde frågan om lämplig rättsliga grund , om den borde vara artikel 37 eller artikel 152 .
jag hänvisar återigen till vad jag sade tidigare om detta och försäkrar henne och kammaren att det skulle vara helt olämpligt för kommissionen att försöka försvara en åtgärd grundad på artikel 37 bara genom att i bestämmelsen undanta varje hänvisning till folkhälsa .
detta är ett ärende som eg-domstolen behandlat vid minst två skilda tillfällen och den har fastlagt rättsliga kriterier för situationer som denna där lämpligheten hos den rättsliga grunden först måste prövas ordentligt när ny lagstiftning läggs fram .
domstolens rättspraxis verkar helt klar med hänsyn till detta .
som en generell kommentar till de här föreslagna ändringarna , särskilt med tanke på frågan om rättslig grund , skulle det vara olämpligt enligt min mening att ändra den rättsliga grunden till artikel 152 under dessa omständigheter då det är mycket troligt att det skulle komma i konflikt med de sakliga kriterier som domstolen lagt fast .
fler av er - nicholson i synnerhet - tog upp frågan om märkning .
i direktiv 70 / 524 förutses frågan om märkning av genetiskt modifierade tillsatser .
det innehåller redan nu texten : &quot; angivelse av särskilda karakteristiska egenskaper på grund av tillverkning av produkter &quot; .
således kommer denna fråga att tas upp .
den formuleringen gjorde det möjligt för oss att ålägga sökanden att i märkningen ange det faktum att genmodifieringsteknik använts i produkten , sakinnehållet i ansökan .
( de ) herr talman ! tillåt mig ytterligare en fråga till kommissionären .
först följande påpekande , kommissionär byrne : europaparlamentet har ingen initiativrätt när det gäller lagstiftningen .
men när ni föreslår en ändring av ett direktiv eller en förordning tar vi oss rätten att titta på hela förordningen och inte bara på den del som ni valt ut .
vi har dessutom i våra ändringsförslag begränsat oss till en formell tillnärmning till andra direktiv . de innehållsliga frågorna har vi till och med avstått från .
de går till exempel inte in på antibiotika .
därför handlar det bara om tillnärmning av de rättsliga bestämmelserna i de enskilda direktiven .
min fråga , kommissionär byrne : vid fn : s konferens i montreal har man just genomdrivit att det i det internationella handelsutbytet måste finnas en märkning av genetiskt modifierade organismer .
tror ni verkligen , att parlamentet - när vi nu har denna möjlighet - kan tillåta att denna märkning inte genomdrivs inom europeiska unionen för fodertillsatser ?
kommissionär byrne , ni är på väg mot en kraftmätning med parlamentet .
vi har förhandlat om lagen om utsäde i två år .
jag ser fram emot våra gemensamma diskussioner .
( en ) jag vill bara understryka att inga genetiskt modifierade organismer har godkänts enligt detta direktiv ; det gäller enbart för tillsatser .
jag vill också säga beträffande frågorna om märkning att detta är en komplicerad fråga .
man håller på att granska detta och skall undersökas på ett allsidigt sätt , särskilt i direktiv 90 / 220 .
denna fråga behandlas just nu av parlamentet och det kommer att bli andra direktiv rörande denna fråga som också kommer att ha artikel 152 som rättslig grund , vilket ger parlamentet fullständig behörighet i fråga om medbeslutande .
jag vill försäkra herr graefe zu baringdorf att det inte alls är min avsikt att få någon sammandrabbning eller styrketest med parlamentet i denna fråga .
min avsikt är som den alltid har varit att samarbeta med parlamentet , att se till att de resultat som vi uppnår är de absolut bästa resultaten .
det bästa sättet att lösa denna fråga är för närvarande genom att lägga fram lagstiftningsförslag för parlamentet , liksom lagstiftningen under utarbetande , snarare än i detta tekniska dokument och under förhållanden där man kanske inte helt har tagit hänsyn till de frågor som läggs fram och som skall diskuteras inom ramen för direktiv 90 / 220 .
det är bäst att avvakta den debatten som enligt vad jag hört skall ske ganska snart .
alla dessa frågor skall tas upp i det lagstiftningsarbetet .
parlamentet noterar era anmärkningar .
skrapie
nästa punkt på föredragningslistan är betänkande ( a5-0023 / 2000 ) av böge för utskottet för jordbruk och landsbygdsutveckling om förslaget till europaparlamentets och rådets direktiv om ändring av rådets direktiv 91 / 68 / eeg i fråga om skrapie ( kom ( 1998 ) 623 - c4-0026 / 1999 - 1998 / 0324 ( cod ) ) .
herr talman , ärade kommissionär ! böges betänkande om åtgärder för bekämpning av tse-sjukdomar hör till de frågor som bygger på de förslag som framförts av parlamentets tillfälliga bse-utskott .
böge har gjort ett betydelsefullt arbete i detta utskott och det är en lättnad att se att det är han som fått i uppdrag att följa upp bse-utskottets arbete i utskottet för jordbruk och landsbygdens utveckling . han har erfarenhet .
jag hade gärna kommit med ett anförande i den diskussionen om man samtidigt hade diskuterat den andra delen av kommissionens förslag .
jag tycker inte det är ändamålsenligt att vi delvis måste föra samma diskussion igen då vi får roth-behrendts betänkande från utskottet för miljö , folkhälsa och konsumentskydd till kammaren .
i föregående inlägg konstaterade schierhuber att skrapie är en mycket förrädisk sjukdom .
för mig som finländare , som har arbetat nära jordbruket i frågor som rör djurens hälsa och transport av djur , är det viktigast att de länder där tse-sjukdomar inte alls förekommer också i fortsättningen garanteras rätten att i tillräcklig grad granska transporter av levande djur .
möjligheten att vid behov granska djuren ytterligare inom dessa områden är inte någon konstgjord protektionism eller någon begränsning av den fria rörligheten när orsaken är välmotiverad .
granskningarna måste ses som rättvisa och kostnadseffektiva handlingar med vilka man främjar djurens välbefinnande och förhindrar att nya kostnader uppstår för eu .
för europeiska liberala , demokratiska reformistiska partiets grupps del kan vi godkänna kommissionens förslag i den mån det gäller böges betänkande , men i behandlingen av nästa betänkande av roth-behrendt måste vi på nytt återgå till situationen i de länder , där tse-sjukdomar inte förekommer .
herr talman ! även jag vill gratulera föredraganden .
det finns inga tvivel om att böge och föredraganden för utskottet för miljö , folkhälsa och konsumentfrågor nu är fantastiska experter på detta område .
det är mycket bra att de fortsätter att bevaka denna fråga på parlamentets vägnar eftersom den är ytterst viktig .
oavsett de många andra angelägna frågor vi har har bse gett oss ett fruktansvärt arv som måste hanteras och lösas .
det är helt klart att förekomsten av skrapie hos får har varit en bidragande orsak till hela problemet .
jag är positiv till den rättsliga grund som läggs fast och till det samlade sättet kommer de nya bestämmelserna hoppas jag att kunna lösa denna situation .
vi måste kunna garantera att ingenting kan införas i livsmedelskedjan eller i djurfoderblandningar så att vi inte låter det som vi tidigare varit med hända på nytt i framtiden .
ingen skulle vilja se att det som hände för bönder med bse någonsin kunde hända igen .
vi måste tillämpa de mest strikta bestämmelser och vi måste få dem att fungera .
det är ytterst viktigt både för producenten och konsumenten att vi återställer förtroendet och det enda sättet vi kan göra det på är genom att ytterst noggrant ta itu med problemet och lösa det .
bse har verkligen inte försvunnit .
man kan hitta det i olika länder .
jag vill inte peka på något speciellt land men många länder står nu inför liknande problem som dem vi hade i förenade kungariket .
den kommer att finnas kvar under ytterligare någon tid .
vi måste se till att hela systemet med spårbarhet och möjligheten att följa djuret från födsel till slakt och rakt genom hela livsmedelskedjan blir en del av den förtroendeskapande mekanismen .
om vi inte kan uppnå det kommer vi att få ofantliga problem i framtiden .
till sist , eftersom jag själv har jordbruksbakgrund har jag under en lång tid absolut trott att om vi hade utfodrat djuren med rätt foder och om djurfodret hade framställts av rätta blandningar skulle vi aldrig haft bse för det första .
det handlade aldrig om bondens ansvar utan det var producenterna av foderblandningar som orsakade detta problem och vi måste försäkra oss om att det aldrig händer igen .
( en ) herr talman ! jag är glad att jag fått detta tillfälle att diskutera en fråga där det finns ett gott samarbete mellan parlamentet och kommissionen , nämligen att bekämpa tse .
jag vill också tacka herr böge för hans arbete i denna fråga .
betydande framsteg har gjorts om vårt förslag till europaparlamentets och rådets förordning om skydd mot och kontroll av tse enligt artikel 152 i fördraget .
detta förslag innehåller alla tse-risker i alla djur och i alla faser i produktionskedjan .
jag är här i dag för att lyssna på era synpunkter på det första steget i denna process för att införa en verkligt omfattande gemenskapssystem för att kontrollera dessa sjukdomar .
i det aktuella förslaget har jag föreslagit att man skall stryka alla nu gällande gemenskapsbestämmelser om skrapie hos får och getter och att införliva dem i ramförslaget om en förordning .
närmare bestämmelser skulle då läggas fram i det ramförslaget .
jag har informerats om att ni är positiva till detta initiativ , vilket verkar vara fallet enligt era bidrag denna eftermiddag , att utforma en enda text .
jag ser fram emot att diskutera varje ytterligare förbättring ni önskar föreslå enligt ramförslaget till lagstiftning , särskilt efter den hänvisning som roth-behrendt gjorde till sitt eget betänkande och ståndpunkt i denna fråga .
jag ser fram emot att få det dokumentet som kommer att beaktas vid alla ytterligare överväganden med hänsyn till denna fråga .
till sist vill jag framföra detta rörande synpunkten att föra in lagstiftningen i bilagor och synpunkten att vi måste uppnå en effektiv balans mellan parlamentets rätt att lämna sina synpunkter och samtidigt vårt krav om snabba resolutioner , snabb lagstiftning och snabba ändringar till gällande lagstiftning .
under de månader jag har varit kommissionär och sett hur lagstiftningsarbetet fungerar i hela systemet inser jag att det krävs mycket arbete på detta område så att vi alla kan uppnå det vi strävar efter , det vill säga överföring av politik till lagstiftning .
gemenskapsåtgärder på vattenpolitikens område
nästa punkt på föredragningslistan är andrabehandlingsrekommendation ( a5-0027 / 2000 ) om rådets gemensamma ståndpunkt ( 9085 / 3 / 1999 - c5-0209 / 1999 - 1997 / 0067 ( cod ) ) inför antagandet av europaparlamentets och rådets direktiv om upprättande av en ram för gemenskapens åtgärder på vattenpolitikens område ) . ( föredragande : marie-noëlle lienemann ) .
( fr ) herr talman , mina damer och herrar kommissionärer , kära kolleger ! vattenfrågan kommer att vara en av de stora miljö- och världsfrågorna under det tjugoförsta århundradet .
om det så handlar om klimatförändringar , världsövergripande resurser , kvaliteten i våra floder och kvaliteten i våra underjordiska vatten , vet vi att de stora utmaningarna medför risker för vår gemensamma framtid .
antingen kommer vi att kunna återställa en vattenkvalitet som motsvarar jordens ekosystem eller så kommer vi att få se en hel rad störningar som hotar utvecklingen i vissa områden och som hotar invånarnas livsvillkor i andra områden , och i grund och botten till och med den globala jämvikten .
som bevis använder jag en utmärkt rapport som vår kollega mario soares har upprättat i de internationella instanserna om havens och oceanernas tillstånd .
när vi talade om klimatförändringar hänvisade vi med rätta till växthuseffekten och atmosfärens tillstånd .
men vi vet också att försämringen av oceanerna i hög grad kommer att destabilisera stora delar av vår jord .
europa bör lämpligen vara så att säga exemplariskt i sina metoder både för att det bör främja en viss modell för utveckling och för att det själv står inför allvarliga problem med föroreningar och vattenförsämring , vare sig det handlar om underjordiska vatten , ytvatten eller hav .
eu har för övrigt undertecknat internationella konventioner . jag tänker särskilt på ospar-konventionen ( international commission for the protection of the north east atlantic ) genom vilken eu har gjort åtaganden .
eu sade &quot; om några år bör vi ha stoppat utsläppen av föroreningar , vi bör ha upphört med att öka föroreningarna och bör till och med närma oss nollstrecket i fråga om giftiga eller farliga ämnen &quot; .
eu undertecknar således de internationella avtalen , därefter följer ett direktiv samt konkreta politiska åtgärder ute i terrängen och då meddelar eu att de fastställda målen inte kommer att kunna uppnås eller också skjuts de upp till sådant datum att själva trovärdigheten i undertecknandet av de internationella avtalen ifrågasätts .
när europaparlamentet tog upp debatten om ramdirektivet om vattenpolitik ansträngde parlamentet sig därför redan vid första behandlingen att kräva en sammanhållning mellan ramdirektivet och de internationella målen samt i synnerhet , när det gäller respekten för ospar , en konvergens som är effektiv och konkret samt stimulerar oss till åtgärder .
eu : s vattenpolitik utgår inte från ingenting .
många direktiv har antagits och kommissionens vilja är för övrigt att lyckas med att göra dem läsbarare , mer överensstämmande sinsemellan samt förse dem med tydligare mål .
det är således en rationell vilja som har lett till genomförandet av detta ramdirektiv .
men parlamentet insisterade vid första behandlingen på att det aktuella direktivet inte bara skall överensstämma med våra åtaganden - typ ospar - utan göra det möjligt för oss att vända på utvecklingen .
för , trots de många direktiven och trots de upprepade förklaringarna om den ansträngning som bör göras i fråga om vattenskydd , när vi ser på miljösituationen i europa , kan vi notera att målsättningarna inte har uppfyllts .
i många fall har situationen förvärrats och vi kan således inte nöja oss med en ansträngning att rationalisera texterna
vi bör sätta upp mål i nivå med de utmaningar som vi har framför oss , och vi har inte mycket tid på oss , för om vi tar för långa frister , såsom kommissionen hade föreslagit , kommer vi inte bara att få ett trovärdighetsproblem hos allmänheten , utan vi vet mycket väl att ansträngningarna kommer att skjutas upp till senare , därefter kommer de att skjutas upp på nytt och således vet man att man inte kommer att nå de uppsatta målen .
jag trycker på denna punkt , för vi får inte vänta oss för hundrade gången att katastrofer rapporteras varje dag i våra tidningar för att säga &quot; jaså ! eu har inte gjort det , jaså !
eu borde ha ... &quot; och då skynda oss att låtsas lösa de problem som man inte ville ta itu med i rättan tid .
exemplet för närvarande med donau och den förorening som sker i rumänien visar mycket tydligt att om vi inte inför en ny ekonomisk utvecklingsmetod , tydliga krav , kontroller och vidtar exakta åtgärder för våra floders tillstånd , vet vi att denna typ av olyckshändelse inte bara kommer att upprepas utan kommer att mångfaldigas med tiden .
vi vet också att om vi inte gör någonting kommer utvecklingen av jordbruket att fortsätta att skapa stor obalans .
floderna i bretagne i mitt eget land är redan nu i en situation av total eutrofiering och det skadar turismen .
herr talman , jag skulle bara vilja avsluta med att säga att det som står på spel är fullt ut klargjort i den andra behandlingen .
vill vi , ja eller nej , ha normer som är förenliga med ospar , det vill säga närma oss noll när det gäller farliga ämnen ?
vill vi förkorta de frister som rådet har föreslagit för detta direktiv ?
vill vi ha en prispolitik som ger möjlighet åt samtliga offentliga och privata aktörer att minska föroreningarna , att verka för föroreningsminskningar och spara vårt vatten ?
vill vi seriöst uppfylla folkens önskningar ?
de flesta ändringsförslag som godkändes av utskottet för miljö , folkhälsa och konsumentfrågor uppfyller denna målsättning , jag hoppas att de kommer att få kammarens stöd .
herr talman , mina damer och herrar ! lienemann har ju nyss redan på ett drastiskt sätt förklarat hur viktigt det är för oss med vatten och luft , framför allt just som grundval för livet för oss människor .
förutom vattenkvaliteten handlar det också om vattenmängden , ty det finns inte heller tillräckligt med vatten överallt i europa , framför allt inte i de mycket torra områdena .
jag beklagar att jag för ögonblicket inte kan se kommissionär wallström här , som egentligen är ansvarig , ty det är hur som helst ett synnerligen viktigt direktiv , som kommissionen har arbetat mycket länge på , och den vattenskyddslagstiftning som vi i dag diskuterar i den andra behandlingen berör alla medborgare i europeiska unionen , men också alla människor i kandidatländerna , som ju måste uppfylla eu : s lagstiftning när de ansluter sig .
vi har arbetat i tio år med denna fråga , och den omfattande ansatsen har blivit möjlig först genom en utfrågning som initierades och genomfördes av utskottet för miljö , folkhälsa och konsumentfrågor .
från den tidpunkten fram till den andra behandlingen i dag har många deltagare i europaparlamentet , kommissionen och ministerrådet arbetat hårt med den .
de 243 ändringsförslagen i utskottet för miljö har vi reducerat till 77 , men nu har ytterligare 30 tillkommit .
ni ser att det finns många frågor , och frågorna är av olika art .
somliga vill ha en skärpning , andra en precisering , många är nationellt präglade .
också i min grupp , europeiska folkpartiets grupp ( kristdemokrater ) och europademokrater , har vi naturligtvis haft olika synpunkter .
vi strävar efter realistiska mål och genomförbara lösningar .
i den andan betyder de ändringsförslag som jag och några kolleger har lagt fram från gruppens sida absolut en förbättring av de krav som föreskrivits i den gemensamma ståndpunkten .
vissa ändringsförslag som vi stöder skall stärka europaparlamentets förhandlingsposition i den kommande förlikningen med ministerrådet .
vi säger klart nej till alla orealistiska krav , som skulle göra europaparlamentet ovederhäftigt .
hit hör för mig nollkravet , dvs. kravet på nollutsläpp fram till år 2020 .
det skulle innebära slutet på all jordbruksverksamhet och mycket av industriverksamheten .
här vill jag än en gång särskilt betona att med de befintliga nationella och europeiska lagarna till skydd för vattnet , hur ofullständiga de än varit och hur litet de än beaktats i medlemsländerna , har vi trots detta redan gjort avsevärda framsteg .
jag vill bara erinra om att vi i dag åter har lax i rhen , vilket för 20 år sedan fortfarande hade varit otänkbart , och att det denna vår skall sättas ut lax till och med i elbe , som varit särskilt förorenad .
det betyder ej att vi inte även i fortsättningen måste göra väldiga ansträngningar för att fortsätta att förbättra skyddet för vattnet och bibehålla den goda vatten- och grundvattenkvalitet som ännu finns , vilket naturligtvis utan tvivel också kommer att vara förbundet med avsevärda kostnader .
många farhågor har just under de senaste dagarna yttrats från jordbrukets sida .
också jordbruk kan bara bedrivas om det finns tillräckligt med friskt vatten till förfogande .
med den linje som vår grupp följt för förhandlingarna med ministerrådet kommer man också att uppnå en bra lösning för jordbruket .
jag bedömer att ledamöterna och allmänheten i detta svåra och delvis mycket tekniska ämne har vilseletts med falska argument från båda sidor .
jag tackar därför i synnerhet mina kolleger i gruppen , som har bidragit med kompromisser .
jag tackar särskilt vår föredragande lienemann för hennes enorma arbete och hennes samarbetsvilliga hållning , även om det fortfarande finns olika uppfattningar på vissa punkter .
men jag tackar också företrädarna för kommissionen , som hela tiden har bistått oss med råd och experthjälp .
om företrädarna för ministerrådet intar en liknande konstruktiv hållning , betvivlar jag inte att vi alla gemensamt kommer att uppnå en ännu bättre lösning för vattenskyddet i europa under förlikningen .
herr talman ! jag vill börja med att gratulera lienemann till det utmärkta arbete som hon har lagt fram och till hennes ansträngningar för att närma våra skilda ståndpunkter i vattenfrågan .
ramdirektivet om vatten är ett nödvändigt initiativ .
om man däremot utgår från att tanken på solidaritet är en reell tanke för processen med det europeiska bygget , är det nödvändigt att man i direktivet tar hänsyn till att vattenresurserna betraktas som en faktor för den sociala sammanhållningen .
vatten - det är det ingen som betvivlar - är en resurs av allmänt intresse .
hanteringen av vattenresurserna förutsätter dock politiska lösningar , när det gäller spanien och andra länder söderut med ett oregelbundet klimat , för att rationalisera förbrukningen samt andra åtgärder för solidaritet .
vi anser att man i detta direktiv bör förespråka en användning av vattnet som gör det möjligt att åtgärda den territoriella obalansen och därför ber jag att ni stödjer ändringsförslag 95 , som har lagts fram av vår grupp .
vi vill säkerställa att artikel 1 i direktivet främjar en hållbar , effektiv , rättvis och solidarisk användning av vattnet .
jag vill nu göra en kort genomgång av de viktigaste punkterna där den spanska socialistiska delegationens uppfattning skiljer sig från de åsikter som försvaras här .
det gäller överföring av vatten mellan magasin .
vi anser att det vore bättre att ett framtida ramdirektiv inte innebar att möjligheten att genomföra dessa är föremål för gemenskapens övervakning .
vi anser med tanke på den spanska statens säregna vattensituation , där överföring sker av strukturell natur , att det bör vara landets myndigheter som beslutar om det egna landets resurser , ett beslut som naturligtvis alltid skall grunda sig på kriterier med sammanhållning och en rationell användning av vattnet som målsättning .
vad beträffar en av de mest omdiskuterade frågorna i vår debatt , nämligen prissättningen , har de spanska socialdemokraterna länge försvarat tanken att direktivet , alltifrån respekten för principen om att &quot; förorenaren betalar &quot; , skall förespråka en policy med rimliga priser på samtliga förbrukningsnivåer .
det är uppenbart att en policy med ett fullständigt återvinnande av vattenkostnaderna inte skulle få samma effekt i spanien som i länderna i centrala och norra europa .
för spanjorerna skulle det innebära att kostnaderna för vattnet ökade för användningen på olika områden , just på grund av de bristande vattenresurserna och för att miljökostnaderna måste inbegripas inom ramen för det som direktivet fastställer .
därför har vi alltid försvarat ett progressivt system för återvinning av kostnaderna , ett system där man har de sociala , miljömässiga och ekonomiska effekterna i åtanke , ett system vars tillämpning anpassas till de olika geografiska och klimatmässiga omständigheterna .
vi vill bygga ett europa med en hållbar och hälsosam omgivning .
men ett miljövänligt europa kan under inga omständigheter byggas i olika hastigheter , utan det bör byggas på en solidarisk grund .
herr talman ! den ekologiska katastrofen i donau påminner oss om hur nära alla länder i europa hör samman och hur viktigt vattnet är för oss alla .
utflödet från kemiska fabriker i min egen valkrets i nordvästra england kommer till slut att hamna på stränderna på europas fastland .
detta klargör de samband som binder oss tillsammans .
detta ramdirektiv är avsett att måla upp en bred skiss för vår politik under de kommande decennierna och det har funnits mycket panik rörande detaljerna .
det är viktigt för oss att komma ihåg att detta är rambestämmelser .
denna skiss är i själva verket mycket generell .
det är lätt för enskilda länder , för enskilda industrisektorer att undkomma de effekter som har målats upp för oss under de senaste dagarna .
det finns många möjligheter att komma undan .
i verkligheten kommer närmare bestämmelser i denna lagstiftning att fastläggas i dotterdirektiv för månader och år framöver .
då är rätta tiden att diskutera några av dessa detaljproblem .
de breda principerna är verkligen sådana som vi borde kunna godkänna - de breda principerna att vi vill minska spridning av riskavfall till grundvattnet , de breda principerna att vi bör inrikta oss på att se till att de kemikalier som vi alla behöver i samhället under alla förhållanden inte bör kunna läcka ut i våra vattensystem .
det finns en kemisk fabrik i nordvästra delen som skrev till mig för att säga att vi måste rösta emot denna lagstiftning .
jag måste fråga dem vad det är för kemikalier som de släpper ut i vattensystemet just nu , och varför de inte meddelar alla som bor i det området exakt vad de håller på med .
detta är något som de helst vill undvika att göra .
principen gäller även vattenhushållning .
den grundläggande insikten som många av oss nu delar är att vi måste införa miljöbeskattning för att uppmuntra till bevarande av resurser , att använda morot och sticka för att få alla att använda våra tillgångar på bästa sätt så att vi inte bidrar till ökad miljöförstöring eller en minskning av en så värdefull resurs som vatten .
jag vill kommentera den politiska positionen här .
den gemensamma ståndpunkten har gjort den ståndpunkt som intogs av parlamentets svagare vid första behandlingen .
några icke-statliga organisationer skulle säga att direktivet i sin nuvarande utformning är sämre än värdelös .
detta är en möjlighet för oss att förbättra situationen .
vi måste vara i stånd att inleda ett medlingsförfarande .
vi har sett omröstning efter omröstning förloras .
åtgärd efter åtgärd har kommit från utskottet för miljö , folkhälsa och konsumentfrågor .
vi har misslyckats med att skapa kvalificerad majoritet .
våra försök att förbättra europas miljö har misslyckats .
vi måste försöka få till stånd ett medlingsförfarande .
vi behöver i slutet av dagen kunna vara säkra på att vi slutligen får en klok och avvägd politik av verkliga förbättringar till rimliga kostnader .
herr talman , kolleger ! redan för nästan trettio år sedan försökte europeiska kommissionen slå fast en europeisk vattenpolitik .
129 kemiska ämnen skulle regleras .
i slutändan fastställdes normer för endast ett tiotal ämnen .
orsaken till det misslyckandet var enhällighetsprincipen .
för ungefär sju år sedan verkade det också som om den europeiska vattenpolitiken skulle offras på subsidiaritetsaltaret .
de konservativa regeringscheferna major och kohl beslutade vid toppmötet i edinburgh att det inte alls var nödvändigt att spanjorer fick lika bra dricksvatten som tyskar och engelsmän .
delvis tränger den inställningen igenom i den gemensamma ståndpunkt som tillkom under det brittiska socialdemokratiska ordförandeskapet .
den ståndpunkten är en ost med hål i , eller för att använda vattentermer , den läcker som ett såll .
det förklarar stormfloden av ändringsförslag från utskottet för miljö : nästan hundra ändringsförslag till den andra behandlingen .
det är ovanligt att göra så men de flesta ändringsförslagen behövs verkligen för att täta alla läckor .
en stor läcka är de farliga kemiska ämnena .
den kemiska industrin och tyvärr även europeiska kommissionen och ministerrådet vill göra en enskild riskanalys för varje farligt ämne .
det tar lång tid , och ännu viktigare , det finns ingen godtagbar nivå för föroreningar genom farliga kemiska ämnen .
endast havets bakgrundsnivå är godtagbar .
det är det som menas med termen &quot; close to zero &quot; .
kommissionen har redan utarbetat en lista med 32 ämnen som prioriteras . många av dessa har en hormonstörande verkan .
det är de så kallade endocrine disrupters . de förorsakar till och med i ytterst minimala mängder könsförändringar hos djur och till och med hos människor , vilket ofta fastställts av vetenskapsmän .
därför är det så viktigt att europaparlamentet uttalar sig för ospar-målet på nästan noll år 2020 .
jag vill ta upp två av de ämnen som finns med på kommissionens lista . kvicksilver och tributyl , förkortat tbt .
på botten av waddenzee ligger värdena för kvicksilver och tbt tio respektive tusen gånger högre än ospar-värdet .
den kemiska industrin och samhället som helhet måste lära sig att byta ut de här farliga ämnena mot oskadliga ersättningar , och om det inte går , att hantera dem i slutna system .
för medlet tbt betyder det att det inte längre får användas som medel för algbekämpning .
mekanisk rengöring av fartygssidorna är ett bra alternativ .
låt mig avsluta med att uttala min förhoppning om att europaparlamentet hämtar upp sin gröna framtoning igen och uttalar sig för nästan noll-alternativet när det gäller farliga kemiska ämnen och hormonstörande ämnen till år 2020 .
herr talman ! i behandlingen av detta direktiv om vatten har parlamentet en avgörande roll .
rådets gemensamma ståndpunkt är helt otillräcklig inom flera områden .
det måste därför nu vara vår uppgift att strama upp och konkretisera kraven i direktivet .
för oss i gue / ngl-gruppen har några principer varit speciellt viktiga när vi har tagit ställning till de olika förslagen .
för det första anser vi att tidsramarna för att genomföra åtgärderna i förslaget måste bli kortare än vad rådet har föreslagit .
vi stöder därför förslagen om snävare tidsramar för att genomföra olika delar av direktivet .
för det andra vill jag att utfasningen av farliga ämnen skall ske på ett konsekvent sätt .
den får inte fördröjas av att man framför nya krav på utvärderingar innan åtgärder vidtas .
i lagstiftningen måste också respekten för internationella konventioner som ospar-konventionen skrivas in .
för det tredje vill vi att prispolitiken skall vara klart uttryckt .
det innebär att grundprincipen måste vara att man betalar de verkliga kostnaderna för vattnet .
i dag får skattebetalarna ofta subventionera industri och jordbruk .
att förorenaren eller förbrukaren betalar skall vara den självklara utgångspunkten för lagstiftningen , även om det också kan krävas undantag i vissa extrema fall .
för det fjärde vill vi att undantagen från reglerna på vattenkvalitetområden skall vara få och tydligt avgränsade .
för det femte vill vi att skyddet av grundvattenkvaliteten och åtgärder mot fortsatta föroreningar i grundvattnet skall vara tydliga och klara .
mot denna bakgrund kan vår grupp rösta för ett flertal av föredragande lienemanns ändringsförslag , såsom de antogs i utskottet .
på ett par punkter skulle vi vilja gå ett steg längre .
vi kommer därför att rösta för de grönas ändringsförslag 102 , 103 och 104 , som vi tycker ytterligare förbättrar positionen .
vad gäller prispolitiken förekommer ibland extremsituationer , som kan kräva undantag från principerna i betänkandet .
jag anser möjligheterna till undantag vara väl tillgodosedda i ändringsförslag 43 från utskottet och uttryckta på ett ännu bättre sätt i ändringsförslag 105 från de gröna .
jag kan inte se att det skulle behövas några ytterligare undantag än de som anges i dessa två ändringsförslag .
detta finns det emellertid olika meningar om inom vår partigrupp .
ändringsförslag 107 , som berör frågan , har lämnats in av en del av vår grupp .
som helhet tycker jag att förslagen från utskottet i lienemanns betänkande är bra , och kan vara en god grund för en svår förlikning .
herr talman ! alla fotografier som tas av satelliter visar att vi verkligen bor på den blå planeten : detta vattenöverflöd är dock en illusion .
den katastrof som nyligen inträffade i donau påminner oss om att floder och älvar är jordens vitala artärer och att föroreningar inte har några gränser .
vatten är en förnybar och begränsad naturresurs .
det minskar då det inte förvaltas på rätt sätt och de geografiska och klimatiska förhållandena inte är gynnsamma .
inom eu är detta en avgörande fråga i medelhavsområdet , men också i andra länder i europa , där vi ser en progressiv uttorkning av våtområden .
känsliga , våta eller torra områden , olikheter mellan stater , olikheter mellan olika regioner inom staterna samt klimatiska , ekonomiska , geografiska , geologiska särdrag är i hög grad bevis som vi vill påminna om men som inte för den skull bör leda till snedvridningar av konkurrensen i gemenskapen .
vi har dock ingett ändringsförslag för att påminna om betydelsen av jordbrukets specifika relation till vatten , en viktig faktor för markanvändning och -bearbetning .
självklart är jordbrukets behov större i söder och detta särdrag måste beaktas i ramdirektivet .
det är för övrigt inte bara i unionens stater som man söker lösningar på dessa problem : partnerskapsländerna i eu-medelhavsområdet begärde i turin i oktober en marshallplan om vatten för medelhavets södra kust .
lyckligtvis är vi inte där ännu .
i europa finns likväl torka , en ökenutbredning av vissa områden , men också översvämningar , och direktivet understryker detta .
vi drabbades nyligen av det i frankrike , också i rhendalen och centraleuropa .
vi behöver detta ramdirektiv såsom en väsentlig beståndsdel av en hållbar utvecklingspolitik , som bör göra de olika användningarna av vatten kompatibla sinsemellan .
men det är nödvändigt att man i denna nya förvaltning införlivar skydd och bevarande av den biologiska mångfalden .
ärendet &quot; vatten &quot; kommer under alla förhållanden inte att avslutas i dag .
frågan om utvidgningen och klimatförändringarna öppnar nämligen nya framtidsutsikter .
herr talman ! vatten av god kvalitet kommer det här seklet kanske att ha ett ännu större strategiskt värde än olja .
det är skäl nog att tacka lienemann för hennes insatser för att ytvattnet skall få en stark ställning .
det verkar vara ganska invecklat att komma fram till en bra ram för den europeiska lagstiftningen .
med ramdirektivet för vattenpolitik vill vi göra slut på den splittrade vattenlagstiftningen i unionen .
därmed undkommer vi emellertid inte ett omfattande och komplicerat direktiv . för det krävs att de verkställande instanserna är mycket noggranna vid genomförandet av det .
särskilt viktigt är det att medlemsstater och vattenmyndigheter utnyttjar sina möjligheter att föra en specifik politik , som tillkommit tack vare tillvägagångssättet med avrinningsområden .
de viktigaste målen förblir att bekämpa en ytterligare nedsmutsning av grund- och ytvattnet , skydda ekosystemen , stimulera en hållbar användning av vatten , bekämpa översvämningar och torka samt att sluta släppa ut farliga ämnen i ytvattnet .
när det gäller utsläppen av farliga ämnen så anser jag att rådets målsättningar är för vaga och inte tillräckligt ambitiösa .
förslaget från miljöutskottet att föra tillbaka utsläppen till nästan noll tycker jag är sympatiskt och eftersträvansvärt .
det måste dock ägnas mycket uppmärksamhet åt genomförbarheten .
därvid måste hänsyn tas till naturliga bakgrundsutsläpp som inte kan påverkas och även svårhanterliga diffusa utsläpp som ändå förorenar vattnet rejält .
herr talman ! vi måste under 2000-talet ta till oss den grundläggande tanken att vi har ett helt nytt förhållande till vattnet .
under 1900-talet var vattnet för oss ett kostnadsfritt transport- och avfallssystem för gift , farligt avfall , kemikalier osv. följderna ser vi redan !
vi måste tänka om och erkänna vattnet som vår viktigaste livspartner , och vårt ansvar för detta går långt utöver de nuvarande generationerna .
på så sätt måste också direktivet behandlas under förlikningen , och befolkningen måste kunna förstå vad vi här planerar , respektive vad kommissionen planerar .
skyddet för vattnet är principiellt också en social fråga , och en avgörande sådan . därför skall principen &quot; förorenaren betalar &quot; användas i större utsträckning , eftersom följderna annars måste bäras av alla .
med tanke på de långtgående skadorna på vattenresurserna är det viktigt att vi inte bara bibehåller nuvarande nivå , utan i morgon vid omröstningen ser till att det skapas verkliga kvalitetsförbättringar .
herr talman ! det är nu redan cirka sex år sedan som vår kollega karl-heinz florenz , assisterad av ursula schleicher , bad om en omstrukturering av hela vattenpolitiken .
det lyckades . det är inget enkelt ämne och jag tycker att de insatser som lienemann gjort förtjänar stor respekt .
beslutsfattandet kring det här ramdirektivet befinner sig i ett mycket viktigt skede .
ämnet har förts in under medbeslutandeförfarandet och vid den första behandlingen har vi därigenom redan kunnat skapa en viktig och sträng lagstiftning .
den gemensamma ståndpunkt som lades fram i slutet av förra året är också en viktig förbättring jämfört med det ursprungliga förslaget .
det är också mycket svårt att föra en politik på den här punkten eftersom skillnaderna är så stora .
till min spanska kollega säger jag : i norra europa har vi ofta översvämningar att tampas med men även förorenat vatten från industrin , medan problemet för kollegerna i söder ofta är att vatten måste transporteras långa avstånd helt enkelt för att ge dricksvatten eller vatten för jordbruket .
jag skall gå in på de två aspekterna av det här ämnet .
först kvaliteten .
nederländerna påverkas till stor del av den europeiska vattenpolitiken .
en mycket stor del , en tredjedel av vårt dricksvatten , utvinns i nederländerna från ytvatten .
nederländerna ligger nedströms , i ett delta , och därför är alltså kvaliteten på det ytvatten som kommer till oss av allra största vikt .
en annan viktig diskussionspunkt är normerna för vattenkvalitet .
i ett antal ändringsförslag sätts det frågetecken för de föreslagna normerna och särskilt med avseende på ospar-normen för år 2020 .
jag förstår väl att vissa tycker att den normen är otydlig eller juridiskt oförsvarlig . jag tycker dock att vi måste stödja den eftersom vi då kan ombesörja noggrannare normer i förlikningsförfarandet .
sedan några ord om kvantitetshanteringen .
en berömd nederländsk poet talade redan i sin dikt &quot; minnen från holland &quot; om vattnet som fruktades på grund av de ständiga katastroferna .
år 1953 inträffade en jättelik vattenkatastrof , varigenom vi samtidigt även blev föregångare när det gäller fördämningar .
år 1990 svämmade våra floder över och vi kunde konstatera att anläggning av konstgjorda verk uppströms påverkar förmågan att ta emot vatten nedströms och kan leda till stora skador .
det betyder att vi även när det gäller kvantitetshantering måste göra stora ansträngningar för att se till att det går bra att leva både uppströms och nedströms .
jag skulle gärna vilja börja med att ge lienemann mina välmenta komplimanger . hon har gjort ett utmärkt arbete .
vatten är ett första livsbehov och en grundläggande rättighet .
var och en borde ha tillgång till rent vatten men tillgång och bra kvalitet på vatten är inte någon självklarhet , det får många erfara , i sydeuropa men nu också i länderna längs donau .
vatten är ofta en källa till konflikter mellan länder och mellan befolkningsgrupper .
därför är det viktigt att vatten blir föremål för internationell samordning .
vi måste erkänna att vatten är vårt gemensamma ansvar .
samarbete inom ett avrinningsområde måste vara en självklarhet .
för liten kapacitet uppströms eller just en för riklig användning kan skapa problem nedströms .
samordning är nyckelordet här .
vattenproblemet blir allt aktuellare .
förändringar i klimatet , små temperaturhöjningar påverkar nederbörden direkt .
vissa områden blir torrare , många områden blir våtare .
i mars anordnas ett andra världsvattenforum i haag .
det här forumet står för en världsomspännande vision .
den visionen måste leda till regionala handlingsplaner för hållbar förvaltning och hantering av vatten .
för europaparlamentet har det nu blivit dags att handla .
vi måste nu ta ställning för en hållbar vattenpolitik som utgångspunkt och samtidigt måste vi vara realistiska .
vi får dock inte heller lägga ribban för lågt .
den gemensamma ståndpunkten är inte tillräckligt ambitiös .
därför är det nödvändigt att vi griper tag i tidigare internationella avtal eller ospar-målen .
vi måste sträva mot en utfasning av farliga ämnen år 2020 .
det är redan avtalat för havsmiljön . det ligger nära till hands att det här avtalet även skall gälla för andra vatten .
ospar-målen håller nu på att utarbetas .
det har ställts upp en lista med 400 ämnen som innebär tydliga risker för miljön .
både tekniskt och ekonomiskt är det genomförbart att i princip minska utsläppet av de här ämnena till noll och det måste vi nu ta ställning för igen .
direktivet skall naturligtvis också vara bindande .
länder nedströms måste kunna lita på att länderna uppströms uppfyller kvalitetsmålen .
kvalitet har ett pris men förorening kan visa sig bli ett mycket högre pris att betala i framtiden .
herr talman , fru kommissionär ! jag vill uttrycka min djupa respekt för det utomordentliga arbete lienemann utfört med detta vattendirektiv .
låt mig påminna om att de riktigt stora miljöproblemen i dag - klimatförändring , skövling av urskogar , utfiskning av haven - hela tiden berör våra gemensamma och absolut nödvändiga , men på något sätt herrelösa resurser .
låt oss också inse att vårt färskvatten i europa kan sägas ligga i gränslandet mellan att ägas av alla och av ingen .
därför är det strategiskt viktigt att ansvaret för vattnet fastställs .
det är också viktigt att de olika vattendragen hålls samman och hanteras som den helhet som de är , oavsett vem som äger den ena eller andra delen av ett gemensamt vattenflöde .
kära kolleger ! förslaget till direktiv utgör i själva verket , som redan flera gånger sagts , en historisk möjlighet att förenkla och förbättra oredan och trasmattan av eu-förordningar och direktiv , och på så sätt uppnå en hög miljöskyddsnivå i europa .
men jag har fått det intrycket att vattenramdirektivets politik präglats av avreglering och åternationalisering .
jag hoppas också att omröstningen inte blir till ett slag i vattnet , och därför är två punkter väsentliga för mig .
för det första ospar .
vi känner till att kommissionens förslag inte går tillräckligt långt ; tyvärr gäller detta också för förslaget från utskottet för miljö , folkhälsa och konsumentfrågor .
att bara slumpmässigt lägga fram förslag , räcker inte .
det vi behöver är ett rättsligt absolut bindande mål för ospar .
endast då kommer vi att kunna åstadkomma rättslig klarhet och framför allt möjligheter till överklaganden .
allt annat skulle förfela sin verkan och inte bidra till att förhindra att ekologiska katastrofer , liknande dem som vi nu upplever i rumänien och ungern , också skulle kunna inträffa hos oss .
jag finner det beklagligt att de nationella regeringarna inte är beredda att engagera sig för ett rättsligt bindande skydd , fastän de ju internationellt har enats om ospar .
men jag tror att det är just det som vi här i parlamentet måste ordna upp , för att därigenom visa att vi inte tillåter att vår trovärdighet utsätts för någon förlust eller någon skada .
det som är viktigt är också att stärka principen om att &quot; förorenaren betalar &quot; , ty priserna måste säga den ekologiska sanningen .
vi får inte ge efter för jordbruks- och kemiindustrins lobbyintressen , utan vi måste propagera och med vår omröstning ge uttryck för att vi vill ha principen &quot; förorenaren betalar &quot; och därmed få kostnadstäckande priser .
vatten är den viktigaste resursen för vårt liv , och vi måste med vår omröstning se till att det finns impulser och påtryckningar för att verkligen iaktta ospar-konventionen .
med hjälp av slutna kretslopp i produktionen är detta möjligt , allt annat skulle vara en urvattning av direktivet .
låt oss ta denna chans !
herr talman ! på den korta tid jag har till mitt förfogande vill jag välkomna föredragandens betänkande och påminna om tre principer som bör vara överordnade de övriga , och som tydligt kommer till uttryck i föredragandens ändringsförslag : vattnet är inte en kommersiell produkt utan något som tillhör unionens folk ; det yttersta målet är att lyckas utplåna alla förorenande ämnen av ytvattnet och grundvattnet , och behovet av att informera befolkningen så att den kan medverka till att återvinna vattnet och inte slösa med det som är en så värdefull resurs .
jag vet att det kan bli problem med det här direktivet , för man talar här om att verkligheten skiljer sig åt i unionens olika länder .
det som händer i norr är inte det samma som det som händer i söder , inte heller som i de länder där man har problem med ökenutbredning .
men vissa ändringsförslag försöker hjälpa länderna i söder , närmare bestämt ändringsförslag 43 som , när det gäller att återvinna kostnaderna , även anger att medlemsstaterna bör ta hänsyn till ländernas sociala och miljömässiga villkor när beslut fattas .
även överledningen av vatten är ett problem .
i mitt land - jag bor i norra spanien - är det stora skillnader mellan norr och söder , och svårigheter uppstår när vattnet skall överledas från en plats till en annan .
men det framgår även av lienemanns betänkande att man i uppsamlingsplatserna bör spara på och värna om vattnet .
jag är medveten om att det är ett komplicerat betänkande , att det finns olikheter beroende på de skilda verkligheterna i länderna , men vi bör föra fram ett ramdirektiv som förhindrar en upprepning av det som händer i donau och det som hände i doñana .
vi kan inte tillåta att man förorenar europas vatten , herr talman , och vi bör upprätta ett direktiv som förstärker regeringarnas politiska vilja att bevara en resurs som vattnet , som är så värdefull för alla .
herr talman ! jag gratulerar föredraganden till ett utmärkt betänkande .
som irländsk ledamot av europaparlamentet som kommer från ett land med stora vattenreserver stöder jag de stora flertalet av förslagen i detta direktiv .
jag skulle emellertid nu vilka granska de sakfrågor som skiljer mellan parlamentets utskott för miljö och rådet .
det senare har redan presenterat sin gemensamma ståndpunkt om denna fråga .
enligt rådet skall målet att uppnå bra ytvattenstatus kunna uppnås senast 16 år efter det att direktivet träder i kraft medan parlamentets utskott för miljö vill få denna tidsfrist förkortad till tio år .
jag ser inget skäl till varför europeiska unionens medlemsstater inte är i stånd att genomföra de centrala bestämmelserna i detta direktiv under så kort tid som möjligt .
jag övergår nu till de ändringsförslag som skall läggas fram för parlamentet i morgon om principen om omkostnadstäckning för vattenutnyttjande .
rådet fastslår i sin gemensamma ståndpunkt att europeiska unionens regeringar måste ta hänsyn till principen om omkostnadstäckning för vattenutnyttjande .
inget bestämt slutdatum för att genomföra denna princip fastslogs i den gemensamma ståndpunkten .
ändringsförslag 43 som innebär att man vill sträva efter att senast år 2010 kunna garantera att vattenprispolitiken i europa skapar tillräckliga incitament för ett effektivt vattenutnyttjande .
vidare skall ett adekvat bidrag från olika ekonomiska sektorer , uppdelat i industri- hushålls- och jordbrukssektorn , garantera att denna politik genomförs .
om dessa ändringsförslag inte stöds i morgon kommer en stark signal sändas ut att mätare och vattenavgifter bör införas för hushåll i alla stater i europeiska unionen .
detta är politiskt opraktiskt ur irländskt perspektiv liksom det faktiskt skulle vara ur andra medlemsstaters perspektiv som portugal , grekland och spanien .
herr talman ! först och främst vill jag gärna tacka lienemann för hennes betänkande .
det är här och nu vi avgör om eu-länderna skall arbeta effektivt för en renare vattenmiljö under de kommande åren .
det gör vi som parlament genom att ändra rådets gemensamma ståndpunkt och visa den väg som leder fram till ett samarbete för en renare miljö .
i oförändrad form kan detta direktiv nämligen få mycket olyckliga och långvariga konsekvenser för miljön och dricksvattnet .
det skulle innebära att man skickade fel signaler till både den europeiska industrin och den europeiska befolkningen .
det är avgörande att stå fast vid en begränsning av det totala utsläppet av kemiska ämnen i våra vattenområden .
det resulterar uppenbarligen i en alltför utdragen tidsaspekt om man skulle göra mätningar av varje enskilt ämne som finns i omlopp , eftersom det finns ca 100 000 .
i detta sammanhang ber jag parlamentet att stödja ändringsförslag 108 , där orden &quot; förorening av vatten genom enskilda förorenande ämnen &quot; , ersatts av &quot; förebyggande av förorening av vatten genom att fortlöpande minska utsläpp &quot; .
vi kan inte försena miljöarbetet genom att överdriva detaljerna i stället för att verka för en minskning av de totala utsläppen av farliga ämnen i miljön .
denna konvention skall vara en riktlinje i arbetet för den rena miljö som vi är skyldiga oss själva och inte minst våra efterkommande .
herr talman ! det är svårt att sammanfatta huvuddragen i ett direktiv som är så viktigt och komplicerat .
i amsterdamfördraget slås fast att vi skall prioritera förebyggande åtgärder , tillämpa principen att &quot; den som förorenar betalar &quot; och skapa en hållbar utveckling där miljökonsekvenserna tas med i beräkningen .
det är viktigt att man urskiljer det ekonomiska värdet av miljöpåverkan vid prissättning och får aktörerna att ta sitt ansvar genom att införa incitament att använda icke förorenande system . detta är odiskutabelt mot bakgrund av förhållandet mellan ekonomisk utveckling och tryggande av miljön , särskilt vattentillgången .
denna situation tar sig specifika uttryck inom många ekonomiska sektorer , men särskilt inom jordbruket .
i det komplicerade förhållandet mellan jordbruk , miljö och vatten , mellan positiva och negativa konsekvenser , mellan en mängd olika lokala situationer och produktionssystem och så vidare , har man infört konceptet om god jordbrukspraxis .
med detta avses den produktionsmetod som används inom jordbruket så att man uppfyller gemenskapens förväntningar på att man skall hålla vården av vattenresurserna på en högre nivå än minimistandarden , med därav följande kostnader och minskade intäkter .
ur detta koncept härrör tvånget att bygga ut och förstärka en integrationsstrategi för att bibehålla vattenvården i centrum av den ekonomiska produktionsmodell som är hållbar mot bakgrund av gällande förutsättningar .
i ljuset av detta skall man inte följa strategin att skilja målsättningen att förhindra att yt- och grundvattnet försämras från målsättningen att skydda , förbättra och återställa dess kvalitet , och därmed skapa en konstgjord prioriteringsskala till förfång för en heltäckande insats med specifika riktade åtgärder inom ramen för denna och där man använder bästa tillgängliga teknik .
vad beträffar att eliminera de föroreningar som härrör från farliga ämnen i vattenmiljön bör man för att optimera tillvägagångssättet införa bestämmelser på både nationell och gemenskapsnivå , så att man bättre kan identifiera de olika typer av vattendrag som förorenats till följd av människors produktion .
slutligen måste man konstruera ett system som innehåller en objektiv förteckning över potentiellt farliga ämnen med mesta möjliga information om kemiska , fysiska och biologiska egenskaper , för att skapa en integrerad modell för insatser på olika strategiska nivåer till skydd för tillgången på vatten som är oundgänglig för oss alla .
herr talman , fru kommissionär , kära kolleger ! om vi tar principen om hållbarhet på allvar , vilken ju är fastslagen i amsterdamfördraget , då kan vårt långsiktiga mål i själva verket bara bli att uppnå nollutsläpp i vårt vatten .
ty vi måste naturligtvis säkra vattnet så att kommande generationer inte belastas av hur vi använder vattnet .
därför gäller det här att utveckla steg med anspråksfulla normer , för att uppnå detta långsiktiga mål . därför stöder jag eftertryckligen lienemanns ändringsförslag för att här utveckla en förnuftig väg med kvalitetsnormer , så att vi verkligen någon gång kan säga att mänsklig användning av vatten faktiskt inte betyder förbrukning av vatten , utan säkrar vattnet i det tillstånd det befinner sig .
direktivet erbjuder några mycket positiva beståndsdelar , som absolut kan framhävas än en gång .
för det första är det den faktiskt breda informationen till allmänheten och delaktigheten för den .
det har det knappast funnits i något europeiskt direktiv .
för det andra är det tvånget till samarbete . jag anser att det är glädjande att man här betraktar vattenresurserna som en helhet och att myndigheter , både i de enskilda medlemsstaterna men också utanför medlemsstaternas gränser , äntligen tvingas samarbeta och se till att det blir en hög nivå på kvaliteten i samtliga vattenresurser .
för det tredje vill jag också ta upp frågan med tidtabellen .
jag är fullständigt övertygad om att vi behöver en strikt tidtabell , så att det också görs ansträngningar för att vi skall nå vårt långsiktiga mål .
jag vill gärna jämföra det med situationen i december .
i december vet vi alla att det är jul den 24 , och vi börjar köpa julklappar .
men hur vore det om vi i december visste att julen skulle inträffa om trettio år ?
vi vet alla hur vi då skulle bete oss . därför behöver vi just när det gäller vattenpolitiken en strikt tidtabell .
jag stöder eftertryckligen föredragandens förslag och anser att vi för alla områden i detta direktiv - vare sig det är en åtgärdslista eller frågan om sysselsättningsåtgärder - behöver en strikt tidtabell .
herr talman ! syftet med detta direktiv bör vara att se till att medlemsstaterna genomför samlade åtgärder för skydd av grund- , dricks- och ytvattnet , och att skyddsnivån motsvarar bestämmelserna i den befintliga gemenskapslagstiftningen på miljöområdet .
låt mig här påminna om att tidigare beslut om nitratdirektivet ännu inte genomförts i samtliga medlemsstater , trots att det är ett gemensamt eu-beslut .
detta förslag innehåller en rad åtstramningar av skyddet för vattenmiljön , som går utöver vårt nuvarande miljömål .
det föreslås att man skall uppfylla ett slutmål för koncentrationer i havsmiljön nära bakgrundsvärdena för naturligt förekommande ämnen och nära noll för syntetiska ämnen skapade av människan .
det är omöjligt och dessutom naturvidrigt .
antagandet av detta betänkande kommer att få allvarliga konsekvenser för jordbruksnäringen i eu , om koncentrationen av t.ex. fosfor och kväve inte får överstiga bakgrundsvärdena för dessa ämnen i vattenmiljön och om man kommer att fastställa ett nollgränsvärde för bekämpningsmedel i vattenmiljön .
jordbruket i europa kommer t.ex. inte att kunna odla brödsäd med förhöjt proteininnehåll , så att säden kan användas till bröd .
resultatet kommer att bli att jordbruksproduktionen flyttar till andra länder utanför eu , med stora sysselsättnings- och samhällsekonomiska kostnader som följd .
jag kan inte rösta för de avsnitt i vattenramdirektivet som behandlar dessa förhållanden .
herr talman , ärade kolleger ! vatten är en dyrbar råvara .
miljoner människor har inte ens tillgång till rent vatten , ett absolut villkor för att överleva .
vi behöver därför inte förundra oss över att vatten ofta är en orsak till krig .
den kapitalistiska världen placerar också ut sina spelpjäser för att få maximal kontroll över vattenförråden .
därvid är det sällan tal om något allmänintresse eller någon solidaritet .
europa står alltså inför en svår uppgift : föra samman den , både när det gäller mål och medel , splittrade vattenpolitiken i gemenskapen i en mer sammanhängande ramlagstiftning .
jag måste bekänna att även i mitt land , flandern , är det en lång väg att gå .
även vi fick nyligen smäll på fingrarna av kommissionen för det .
varje förnuftig människa vill att det här ramdirektivet används som ett påtryckningsmedel för de politiska ledare som nu kommer till korta .
den gemensamma ståndpunkten är i det avseendet en fars , ett verk utan tvång , en riktig förolämpning mot ospar-avtalen .
vi har till och med en tidsfrist för genomförande som kan tänjas ut till 34 år framåt .
mina barn kommer då att vara äldre än vad jag är nu .
håll med om att det här inte är rätt .
i morgon kan vi välja en svag ram utan tvångsmekanism som förgiftar framtiden för våra barn .
antingen röstar vi för ändringsförslagen från min grupp , från föredraganden eller från utskottet för miljö .
de senaste månaderna har det varit en enorm lobbyverksamhet på gång .
vad som var iögonenfallande i den här saken var den enorma pressen från ministerrådet .
i mitt eget land skedde det både genom de flamländska och de wallonska miljömyndigheterna .
de ställer sig bakom den svaga gemensamma ståndpunkten till förmån för ett ytterligare ställningstagande av vårt parlament .
jag undrar verkligen om det här är ett försök som de gröna miljöministrarna i mitt land känner till .
kolleger ! det räcker inte längre med vackra ord .
vi måste göra en resolut kursändring .
vid omröstningen i morgon kan vi göra det tydligt att europa anstränger sig för att skapa en ansvarsfull och framtidsinriktad vattenpolitik .
det kan bara öka vår trovärdighet .
jag förklarar debatten avbruten och den kommer att återupptas kl. 09.00 .
dialog om europa : institutionella reformens insatser
nästa punkt på dagordningen är kommissionens meddelande - dialog om europa - institutionella reformens insatser .
i kommissionen pågår just nu en debatt och mycket skall till för att detta arbete skall avslutas i dag .
jag kommer huvudsakligen för att , såsom angetts på föredragningslistan , tala om ett nytt initiativ som kommissionen förslår till svar , och det är inte det enda svaret , på en stor utmaning som bör mobilisera samtliga aktörer i den europeiska uppbyggnaden , i vilken ni befinner er i första ledet i egenskap av parlamentsledamöter , men också jag såsom kommissionsledamot , också de ministrar som sitter i rådet , de nationella parlamentsledamöterna och jag vill tillägga till och med de tjänstemän som arbetar i de olika institutionerna och som är engagerade i och motiverade av denna europeiska uppbyggnad .
i den långa debatten i morse där jag deltog vid sidan om ordförande prodi berörde många av er det demokratiska underskottet och det stora avståndet till de europeiska institutionerna .
när jag säger det försöker jag inte bara att ställa frågan - en av er sade det mycket tydligt och med stor kraft : vem gör vad ?
och det minsta man kan begära är att medborgarna förstår vem som gör vad i våra olika institutioner .
frågan ställs då omedelbart också om vad vi gör tillsammans och vad vill vi göra tillsammans i framtiden , i synnerhet med de länder som skall ansluta sig till oss .
det demokratiska underskottet får oss således också att undra och därför beslutade vi nyss i kommissionen att redan dagen efter öppnandet av regeringskonferensen , under vilken jag har fått äran att företräda kommissionen vid prodis sida , och i nära samarbete med era båda företrädare , brok och tsatsos , lägga fram &quot; en dialog för europa och om europa &quot; och att för vår del delta i direktkontakten med medborgarna .
samtliga kommissionsledamöter har åtagit sig att varje gång som de måste bege sig till ett land , och inte bara sitt ursprungsland , och till ett område - för min del händer det tre eller fyra gånger per månad - ägna ett ögonblick av sin tid åt en direktdialog med medborgarna , inte bara med eliten eller de institutionsansvariga som man vanligen möter utan också skapa en direktkontakt i ett universitet , ett gymnasium eller en fabrik , att söka kontakt med människor , svara på frågor och lyssna .
det kommer att bli den del som vi tar på oss , såsom ni kommer att göra det själva när det gäller denna nödvändiga ansträngning och angelägna förpliktelse som består i att minska det demokratiska underskottet , det vill säga avståndet till medborgarna i förhållande till vad vi gör .
vi vill att detta initiativ skall skötas i samarbete med medlemsstaterna och i förbindelse med europaparlamentet .
vi kommer att göra en regelbunden sammanfattning så att den allmänna opinionen mäts och man kan justera eller omorientera .
vi vill också agera i samråd med de nationella parlamenten , de lokalt folkvalda , icke-statliga organisationer , arbetsmarknadens parter och media .
opinionsnätverk , politiska grupper och partier , europaparlamentets ledamöter , nationella parlamentsledamöter , folkvalda , det sade jag just lokala myndigheter eller nationella parlament , regionkommittén , ekonomiska och sociala kommittén , det civila samhällets organisationer och universitetsmiljöerna kommer att beröras .
jag vill för övrigt påminna om - behöver jag göra det - att europaparlamentet själv redan tog initiativet den 1 februari , och jag vill åter tacka ordförande napolitano för det , att ordna ett första arbetssammanträde med företrädarna för de nationella parlamenten , det vill säga företrädare för medborgarna i varje stat .
kommissionen kommer att föreslå medlemsstaterna att ansluta sig till denna åtgärd , antingen inom ramen för ett tillfälligt samarbete eller i ett mer strukturerat partnerskap .
vi upprättar en plan för media och nära kontakter med eu : s ordförande och europaparlamentets talman .
jag har sagt på vilket sätt kommissionsledamöterna kommer att delta vid möten och besök ute bland människor .
vi vill ha medborgardebatter .
kan jag bara , utan att föreläsa - framför allt inte - och inte heller ge råd , påminna om att när jag hade äran att vara minister för europafrågor i mitt eget land , kände jag behovet av att få en direktdialog med medborgarna och när jag varje vecka förde den dialogen direkt i olika områden upptäckte jag att det fanns ett enormt behov av att ge ett ansikte åt europeiska unionen och jag åkte således med en ledamot från europeiska kommissionen , inte bara de franska kommissionsledamöterna för övrigt , ambassadörer i tjänst i paris , ledamöter från europaparlamentet , och förde en dialog och jag upptäckte att det fanns oändliga frågor , att de var intelligenta , att människorna hade ett behov av att respekteras , att man lyssnade till dem och förklarade för dem .
det är vad vi skall göra med stöd av ett budgetanslag på omkring fyra miljoner euro som vi ber er ställa till vårt förfogande .
det kommer att bli nödvändigt att förhandla fram ett anslag inom ramen för budgeten år 2001 för vi vill föra fram och leda denna idé inte bara försöksmässigt , utan varaktigt år 2000 och 2001 , det vill säga under hela förhandlingen i regeringskonferensen och ratificeringsprocessen .
vi kommer att inleda denna dialog i bryssel den 8 mars i närvaro av sjuhundra unga provanställda i kommissionen .
er talman , nicole fontaine , har accepterat att stå vid ordförande prodis och flera kommissionsledamöters sida för att inleda den första dialogen och , mina damer och herrar ledamöter , jag kommer att se till att varje gång en kommissionsledamot inleder en dialog skall de ledamöter från europaparlamentet som finns närmast tillgängliga kunna vara närvarande själva och ge sin synpunkt och förklara europaparlamentets arbete och roll .
ja , det var vad jag ville säga , herr talman .
jag är för övrigt beredd att svara på frågor , ta emot idéer och förslag från de ledamöter som är här .
kolleger , ni känner till bestämmelserna .
ni förväntas ställa frågor och inte nödvändigtvis göra långa uttalanden .
ni har en minut var att ställa er fråga .
herr talman ! jag vill ge uttryck för min och , tror jag mig kunna säga , utskottets för konstitutionella frågor , vars ordförande jag är , uppskattning av detta initiativ från kommissionen .
detta initiativ motsvarar för övrigt de anvisningar parlamentet självt gav i sin resolution från den 18 november .
jag har också hört de preciseringar kommissionär barnier gav om förhållandet med och kopplingen till europaparlamentet när detta program utformades .
om ni tillåter kommissionär barnier , skulle man inte i meddelandetexten kunna säga någonting mer om detta än den enkla , litet kalla , frasen &quot; elle sera conduite en liaison avec le parlement européen &quot; ?
jag tycker att det vore bra om man kunde betona denna överensstämmelse i avsikter och bemödanden , även eftersom jag kan urskilja ett speciellt samordningsproblem som är just det mellan kommissionens initiativ , som verkligen inte bara riktar sig till ledamöter i europaparlamentet utan även till ledamöter i nationella parlament och vårt utskotts program .
efter den studiedag den 1 februari som kommissionär barnier hänvisade till och där kommissionens betydande bidrag var till stor nytta är vår avsikt att ta upp regeringskonferensens utveckling vid alla våra möten .
vi kommer därför att ha ledamöter i de nationella parlamenten närvarande vid alla våra möten , ett kvalificerat och bestående deltagande hoppas vi , och detta kommer att bli en kanal som blir ett bra komplement till dem i kommissionens initiativ .
tack , ordförande napolitano , jag bekräftar att det vi föreslår överensstämmer fullt ut med andan i resolutionen av den 18 november och jag vill också här säga att jag har kunnat föreslå kommissionen detta initiativ tack vare min kollega vivianne redings samarbete och goda samförstånd samt att det genomförs i förbindelse med günther verheugen , eftersom allt som står på spel och de stora utmaningarna , som vi måste förklara och våra landsmän i varje land undrar över och frågar om , gäller både utvidgningen - utvidgningens möjligheter och risker - och den institutionella reformen .
jag har mycket väl förstått er oro , ordförande napolitano , och det kommer att bildas en interinstitutionell arbetsgrupp ( det första sammanträdet kommer att äga rum i mars ) .
jag skall se till att vi går bortom det som litet torrt står i kommissionens text , att vi talar om mer än förbindelse , om gemensamt arbete och att man sålunda under dessa två år kan samordna de initiativ som ni tar och som vi tar , var och en å sin sida , men som vi tar tillsammans .
mina damer och herrar ledamöter , låt mig säga att om vi vill inleda denna dialog finns det arbete för alla .
herr talman , herr kommissionär ! det är ljuv musik för mina öron att höra er nämna ordet medborgare så ofta .
i detta parlament talar man mer och mer om den allmänna opinionen : rädsla för allmänna opinionen , det är som ni vet litet paternalistiskt , men vårt parlament är nu en gång så och vi måste acceptera det .
jag ville ställa en exakt fråga till er inom ramen för frågan om regeringskonferensen : jag tror mig veta att domstolen i luxemburg håller på att noggrant behandla en viktig fråga som handlar om bedrägeribekämpning och olaf .
såsom ni vet finns det förvisso problem som berör parlamentet men också europeiska tjänstemän , för de är också europeiska medborgare .
jag ville fråga er med tanke på hur brådskande denna fråga har blivit om kommissionen har tänkt på möjligheten att ändra struktureringen av organisationen för bedrägeribekämpning fullt ut genom att tänka ut en lösning som innebär att bedrägeribekämpning i medlemsstaterna liksom i de europeiska institutionerna skulle ingå i domstolens behörighetsområde .
herr dupuis , först och främst sätter jag stort värde på ordet medborgare i mitt offentliga liv .
det är ett av de finaste orden i en demokrati och jag tror att det måste användas .
vi skall föra en dialog med medborgarna , inbegripet med de anspråkslösaste eller med de människor som är längst bort ifrån besluts- och informationscentrerna .
eftersom ni talar om regeringskonferensen vill jag bara med anledning av frågan om bedrägeribekämpning i synnerhet - om det nu handlar om att kämpa mot bedrägeri mot gemenskapens intressen och budget - påminna om att vi för övrigt i kammarens arbetsanda och kanske genom att gå samma väg , kan jag säga att vi tagit fasta på idén i kommissionens förslag om att inrätta en speciell och ny tjänst såsom europeisk åklagare ; denne skulle således ha befogenhet enligt fördraget , således av medlemsstaterna , att från början till slut undersöka ett ärende som eventuellt ifrågasätter gemenskapens intressen och budget .
vi noterar helt klart och nästan kliniskt att det rättsliga samarbetet inte längre räcker till , inte räcker för närvarande för att effektivt kunna bekämpa dessa bedrägerier , var de än kommer ifrån , inifrån eller utifrån , och därför har vi lagt fram detta förslag om att inrätta tjänsten som europeisk åklagare , som efter att själv ha undersökt ett ärende från början till slut skulle kunna låta det undersökas därefter och dömas av lämpligaste nationella domstol .
vi har inte - jag svarar på den andra punkten om domstolen - vi har ännu inte klargjort våra ståndpunkter om domstolen eftersom vi väntade på betänkandet dur som inlämnades för några dagar sedan .
såsom jag hade åtagit mig skall kommissionen komplettera sina förslag rörande yttrandet om regeringskonferensen , i fråga om domstolssystemet och domstolen , inom de närmaste veckorna .
herr talman , herr kommissionär ! i förrgår visades en toppnyhet i det mest sedda danska nyhetsprogrammet , som jag vill be er kommentera .
historien handlade om att en tjänsteman i kommissionen skulle ha sagt till en företrädare för det österrikiska näringslivet att eftersom han var österrikare så kanske han skulle utestängas från deltagande i ett vetenskapligt utbytesprojekt tillsammans med företag i andra länder , inklusive danmark .
jag vill be er att bekräfta att om en tjänsteman har sagt att ett österrikiskt företag på något sätt skall utestängas från deltagande i gemensamma utbytesprojekt , så har denna tjänsteman uttalat sig på ett felaktigt sätt , och om han inte har sagt så finns det ingen historia .
herr haarder ! enligt min vetskap har ingen tjänsteman fått tillstånd att säga något liknande .
det skulle inte vara , här uttrycker jag min personliga åsikt , normalt och rättvist att straffa de österrikiska medborgarna , företagen och de anställda på grund av oro över att en ny koalitionsregering bildats i detta land .
med reservation för en kontroll som jag skall göra eller låta göra omedelbart efter sammanträdet bekräftar jag således vad jag sade : kommissionen har aldrig sagt eller beviljat något i den stilen .
herr haarder , det finns annat som vi rent allmänt kan lära oss av det som händer i österrike .
jag har själv tagit upp olika möjliga svar på denna utmaning som för oss alla består i att påminna om och att på nytt visa vad vi gör tillsammans sedan 1957 : en ekonomisk gemenskap , naturligtvis , men först och främst en värdegemenskap och en stadga om grundläggande rättigheter som kommer att mer och tydligare skydda enskilda medborgare , artikel 13 i fördraget rörande diskrimineringar .
vi föreslog redan före den österrikiska krisen i vårt yttrande av den 26 januari att denna artikel efter regeringskonferensen skall omfattas av kvalificerad majoritet och inte längre av enhällighet , och det finns en eventuell möjlighet , jag säger eventuell , - det säger jag personligen - att komplettera artikel 7 med en ny strecksats som skulle förse förfarandet med övervakning eller demokratiskt larm på rättslig grund och sedan slutligen offentlig debatt .
det enda sättet att få bort dåliga idéer är att ersätta dem med nya .
jag återvänder därmed till ämnet för diskussionen : just nu tror jag djupt på debattens demokratiska värde och kraft , i synnerhet för att bekämpa demagogi .
kommissionär barnier ! ni lade stor vikt i er redogörelse vid hur viktigt det är med en dialog med europas medborgare .
med hänvisning till regeringskonferensen , som ni vet , tilldelades enligt besluten i helsingfors det portugisiska ordförandeskapet en speciell rätt att utöka dagordningen för konferensen under konferensens gång .
utan tvivel har parlamentet sina egna företrädare , brok och tsatsos , närvarande .
men kan ni , herr kommissionär , även lämna ett löfte att om och när dagordningen utökas av rådet så skall ni meddela detta till parlamentet så att vi kan diskutera det mellan oss själva och naturligtvis med er med avsikten att fortsätta den dialogen med medborgarna som ni lagt så stor vikt vid ?
( fr ) herr beazley ! mitt svar är ett klart och tydligt ja , men det är uppriktigt sagt ingen nyhet .
ordförande napolitano , många ledamöter från utskottet för konstitutionella frågor och ännu fler ledamöter här i plenarsammanträdet vet att jag kommer att vara tillgänglig för att under hela förhandlingen på kommissionens vägnar tala om hur det går i en anda av öppenhet och på realtid .
jag kommer kanske att säga det på annat sätt än professor tsatsos och elmar brok som är era direkta företrädare . det är för övrigt troligt att vi kommer att säga det tillsammans vid många tillfällen .
jag tror att det är viktigt att förhandlingen inte är hemlig vare sig för europaparlamentet eller för de nationella parlamenten , vilka , vill jag påminna om , i sista hand måste avge sin åsikt och inta en ståndpunkt i ratificeringsprocessen .
därför hyllade jag napolitanos initiativ till ett gemensamt och regelbundet samråd mellan de femton ländernas nationella parlament och europaparlamentet .
därmed börjar öppenhets- och debattskyldigheten här när det gäller institutionsreformen .
jag kommer således att vara tillgänglig varje gång ni önskar det för att redogöra för våra ståndpunkter och framstegen i förhandlingen under hela detta år .
herr talman ! i första hand mina komplimanger för kommissionens handlingssätt .
jag tror att det är mycket bra att man inleder samtal med medborgarna i ett tidigt skede , det skedde ju inte vid amsterdamfördraget eller vid maastrichtfördraget och det har bara lett till en stor misstro .
två frågor : för det första , ni har sagt att ni skall samtala med medborgarna och jag börjar redan med 700 praktikanter vid europeiska kommissionen .
tänker ni också rikta er till medborgarna via media , alltså även via tv och via internet ?
min andra fråga är en kritisk fråga .
det har nyss lagts fram ett förslag om öppenhet och insyn från europeiska kommissionen .
om jag jämför det med det förslag som gäller för lagstiftning hos oss i nederländerna så är det bara en liten skugga av det och det förslaget har lett till mycket kritik i nederländerna .
min fråga är egentligen : hur vill ni utforma öppenheten med avseende på regeringskonferensen , det direktiv som nu lagts fram är nämligen inte något bra exempel på det .
fru ledamot , fru minister maij-weggen , eftersom vi talar om öppenhet när det gäller regeringskonferensen vet ni hur det kommer att gå till . förhandlingen börjar för övrigt just i detta ögonblick .
representantgrupperna har sammanträde i bryssel och jag skall skynda mig till dem strax .
dokumenten kommer för det mesta att vara öppna , arbetsdokument .
vi kommer inte att diskutera inför media under förhandlingssammanträdena som kommer att pågå under hela året mellan ministrarna och europeiska rådet men jag har åtagit mig , jag kan inte göra annat just nu , att genomföra denna öppenhet och att redovisa i institutionerna om förhandlingen och om kommissionens ståndpunkt .
jag vill bekräfta , samtidigt som jag tackar er för att ni frågat mig om det , att vi kommer att använda alla moderna medel , i synnerhet television , för att sända de offentliga debatterna i det ena eller andra landet , och till och med på europeisk nivå .
vi kommer att öppna ett forum på internet och skapa permanenta fora för diskussioner .
kommissionsledamöterna skall åta sig att snabbt svara på alla frågor som ställs .
vi kommer att använda alla dessa moderna medel .
men jag tror att vi också måste anstränga oss att gå så nära inpå människorna som möjligt .
jag skulle vilja att i samtliga europas regioner - det är utan tvivel ännu litet utopiskt - skall en kommissionsledamot , när han kan det , en ledamot från europaparlamentet , eller en minister kunna gå till offentliga debatter .
jag har bevis för att det är möjligt .
de flesta av er gör dessa debatter i era valområden och i era regioner .
ur kommissionens mer egoistiska synpunkt skulle jag vilja att denna institution får ett ansikte i medborgarnas sinnen och att de män och kvinnor som utgör den skall så ofta som möjligt kunna gå medborgarna till mötes .
herr talman ! jag uppskattar barniers löfte att gå ut till regionerna , både för att förklara och för att lyssna till vad medborgarna har att säga .
jag skulle vilja inbjuda honom till min egen region , yorkshire , en större europeisk region som är en fullvärdig deltagare på den europeiska inre marknaden och en mycket stor mottagare av europeiska strukturfonder .
han kan komma med båda de hattar han bär som en kommissionär .
jag skulle vilja fråga honom hur energiskt kommissionen kommer att satsa på denna informationskampanj ?
i några medlemsstater är det inte bara fråga om att tillhandahålla information till en allmänhet som inte är så välinformerad som den kunde vara .
det är naturligtvis viktigt men det gäller också att bekämpa den felaktiga information som sprids av en mycket aktiv anti-europeisk rörelse och av de anti-europeiska organisationer som finns .
kommissionen måste ge mycket kraftfulla svar på några av de synpunkter som den kommer att få ta emot som en del av kampanjen .
herr corbett , jag tackar er för er uppskattning .
jag accepterar gärna er inbjudan och om jag har förstått rätt , vill ni att jag , när jag kommer till yorkshire , inte bara tar upp reformen av de europeiska institutionerna utan också strukturfonderna .
jag kommer således att besöka er för att genomföra denna dubbla uppgift .
jag glömde för övrigt att tala om hur angelägen jag är att möta , och jag har redan gjort det , de nationella parlamenten , inte bara genom att träffa deras företrädare här , utan genom att åka och träffa dem på plats .
för tio dagar sedan var jag i westminster . ni ser , herr corbett , att jag inte är rädd för svårigheter .
jag skall nästa vecka besöka bundestag i berlin .
jag har varit inför den franska senaten .
under hela denna debatt kommer jag således att också varje gång det är möjligt direkt besöka de nationella parlamenten .
vad beträffar dialogen med medborgarna handlar det inte om att göra propaganda eller marknadsföring , inte ens kommunikation .
jag skulle vilja att dialogen verkligen blir en dialog , och att efter en liten film som objektivt förklarar vad som står på spel i fråga om den institutionella reformen , skall de som är här på tribunen kunna uttala sig och svara direkt .
vi skall , jag upprepar det , genomföra detta initiativ till dialog i tillfälligt eller strukturerat samarbete med medlemsstaterna och jag vill mycket gärna med ert stöd att de femton medlemsstaternas regeringar skall kunna ansluta sig på de sätt som de anser lämpliga och passande till detta initiativ till dialog .
herr talman ! jag vill gärna ansluta mig till barniers diskussionsgrupp med de 700 provkandidaterna , så han har några att diskutera med .
det är ju inte så roligt att bara diskutera regeringskonferens och öppenhet med sig själv .
under framställningen i parlamentet sade barnier , i samband med regeringskonferensen , att socialpolitiken inte var underställd majoritetsbeslut , men när jag tittar på sidan 63 ser jag att kampen mot olika behandling , rätten att resa och att bosätta sig - alltså bosättningsdirektiven - hela socialförsäkringen , förnyelsen av förordning 1408 , av åtgärder på det socialpolitiska området - med ett fåtal undantag - skall underställas majoritetsbeslut .
förstår inte barnier att han går inte i hjärtat av medlemsstaternas valförfaranden ?
det är ju p.g.a. dessa frågor som folk går till val och som leder fram till en ny majoritet i folketing och andra parlament .
kan det styras från bryssel ?
är det ett led i den genomgripande decentralisering som prodi talade om i förmiddags ?
jag blev mycket glad när jag hörde förra veckan att kommissionen under flera år noga skall granska begreppet subsidiaritet avseende inte bara förbindelserna mellan union och medlemsstater utan också union , medlemsstater , regioner och städer .
jag hoppas att kommissionär barnier i sin strävan efter dialog i europas regioner kommer att utveckla den tanken och lära av det han får höra .
jag hänvisar till ett av era svar på de föregående frågorna där ni nämner det som jag kallar låsningen av fördraget inför snedvridningsriskerna , i synnerhet den mångfalden av sanktioner som kan drabba en medlemsstat genom tillämpning av artikel 7 för brott mot grundläggande fri- och rättigheter .
tror ni att dessa förslag , eller förslag av denna typ , kan ingå i regeringskonferensens uppgift såsom den definierades i helsingfors ?
jag har för min del inte det intrycket .
är ni inte rädd för att sådana sanktioner skall kunna slå slint och användas till att straffa , inte brott mot mänskliga rättigheter , utan små skiljaktigheter , åsiktsförbrytelser eller åsiktsskillnader i förhållande till den dominerande europeiska tanken ?
ja , herr bonde , vi kommer att inleda debatten med sjuhundra ungdomar i bryssel .
det är så att de kommer att arbeta i institutionerna och hos kommissionen och jag tror att det är bra att inleda debatten med ungdomar som är motiverade .
när det gäller det sociala trygghetssystemet vill jag bekräfta att vi har lagt fram förslag på området för kvalificerad majoritet eller på området för enhällighet utan ideologi .
i ert land , bonde , liksom överallt tror jag att man är angelägen om att den inre marknaden skall fungera bra på de mest rättvisa villkor för konkurrens och rörlighet för varor och personer .
och det är således det som är vår regel .
vi föreslår nämligen att vi skall besluta med kvalificerad majoritet om vissa politiska områden , vissa skatteåtgärder eller i fråga om social trygghet och hälsovård när det har ett direkt samband med den inre marknadens funktion .
vårt förslag är inte övergripande och det är inte systematiskt .
jag känner mycket väl till hur känsliga dessa frågor är om beskattning och social trygghet .
jag tror inte att vi skall stöpa samtliga nationella system för social trygghet i samma form , det har aldrig varit fråga om det , utan helt enkelt att säkra bästa villkor för den inre marknadens funktion i ett europa med trettio eller tjugosju länder utan att en stat skall kunna låsa de tjugosex eller tjugosju övriga staterna .
herr maccormick , ja , jag bekräftar att denna dialog bör gå utanför de nationella huvudstäderna och att den bör gå så nära inpå människorna som möjligt , där de bor och har sina rötter och om jag sade något annat skulle jag inte vara överens med mig själv i egenskap av kommissionär med ansvar för regionalpolitik , det vill säga ett av de konkretaste och synligaste politikområdena , som är gjort för att stödja sysselsättning och livskvalitet för människor i regionen och ni kommer ofta att få höra mig säga att denna politik inte bara har skapats för det prioriterade målet med sammanhållning och solidaritet mellan regionerna , den har också skapats såsom ett komplement för att människorna skall kunna behålla sina rötter , sina traditioner , sin själ och sin identitet där de bor .
vi skall således föra denna dialog med städer och regioner .
berthu , helsingforsmandatet är klart och tydligt och vi är inom denna ram .
där planeras att de tre grundläggande ämnena som åsidosattes i amsterdam skall behandlas först och prioriteras .
tillhörande institutionella frågor läggs till samt slutligen frågor som det kan bli lämpligt , beroende på de portugisiska och franska ordförandeskapen , att tillföra under förhandlingen .
kommissionen spelar sin roll om den tror att den bör komplettera i den ena eller andra frågan sitt yttrande som behandlar många institutionella frågor .
jag är ännu inte säker på att vi kommer att göra det om artikel 7 och om vi gör det kommer vi inte bara att göra det till svar eller reaktion på en konjunktursituation , som är tillräckligt allvarlig för att de fjorton regeringarna i unionen har mobiliserats tillsammans för att lämna sitt svar och vi kommer också att göra det med tanke på framtiden i allmänhet .
alla medel som definitivt kan stärka den värdegemenskap som vi utgör tillsammans alltsedan unionen grundades 1957 och till och med tidigare på ruinerna av andra världskriget , allt som kan göras kommer att vara lämpligt .
herr berthu , jag är säker på att vi kommer att kunna bli överens , ni och jag , på denna grund .
ni har besvarat frågorna noga och även inlett den dialog om europa som hänvisade till .
ni har visat ett mycket gott exempel på hur man håller tiden i dag .
det avslutar debatten .
nästa punkt på föredragningslistan är frågor till kommissionen ( b5-0009 / 2000 ) .
fråga nr 36 från ( h-0025 / 00 ) :
angående : hög barnadödlighet i kosovo enligt världshälsoorganisationens senaste uppgifter till fn har kosovo högst barnadödlighet i europa ; nästan 50 procent av alla för tidigt födda barn dör . till följd av kriget har missfallen ökat kraftigt och de barn som inte föds för tidigt är mindre utvecklade än normalt .
kan kommissionen , mot bakgrund av den humanitära hjälp som eu tillhandahåller och det politiska sändebudet bernard koushners ansträngningar , meddela vilka åtgärder den har vidtagit till skydd för kvinnorna i kosovos rätt till moderskap och för gravida och födande kvinnors samt spädbarns hälsa ?
herr talman ! kommissionen är medveten om den mycket svåra situationen i fråga om hälsovård och hälsovårdsanordningar i kosovo , inte bara för gravida kvinnor utan på hela fältet .
detta beror både på den senaste konflikten och på alla år före konflikten av misskötsel och brist på underhåll .
den statistik som nämns i fråga om barndödlighet talar för sig och är helt oacceptabel .
situationen är dock knappast bättre för andra delar av befolkningen .
kommissionens svar har varit följande : först och främst har hälsosektorn fått motta betydande bidrag från echo .
echo inriktar sig för närvarande på att tillhandahålla medicinsk utrustning och akut hälsovård , på stöd till inrättningar liksom vaccinering .
insatserna inriktas dock alltmer på att upprätta ett självförsörjande hälsovårdssystem i provinsen .
unmik har redan tagit på sig en betydande roll på detta område .
vidare har det i enlighet med återuppbyggnadsprogrammet inletts brådskande insatser på sjukhuset i mitrovica i form av ett återuppbyggnadsprogram på 1 miljon euro .
utvecklingen går långsamt på grund av de spända förbindelserna mellan de etniska grupperna i denna delade stad .
kommissionen fortsätter dock sina insatser med stöd av unmik för detta projekt .
vi hoppas att det en dag blir en symbol för att främja fördelarna med etnisk försoning .
enligt europeiska gemenskapens uppskattning av skador uppgår de beräknade kostnaderna för återuppbyggnad av hälsovårdsinrättningar och anskaffning av utrustning till apotek och vårdcentraler till 4 miljoner euro .
kommissionen skall nu inleda arbetet med biståndsprogrammen för år 2000 .
vi tror att vi kan anslå en betydande summa till att förbättra hälsovårdssystemet .
tonvikten kommer att ligga på långsiktiga reformer som täcker finansiering liksom utbildning och materialanskaffning inom hälsosektorn .
arbete pågår redan tillsammans med unmik för att fastslå ett lämpligt bidrag från kommissionen för detta initiativ .
herr kommissionär ! i morse framhöll ordförande prodi bl.a. att vår förmåga till effektiva insatser sätts på prov på balkan , att europeiska unionens trovärdighet sätts på prov och att det är dags att låta ord och handling följas åt .
vi har fått uppgifter om den höga spädbarnsdödligheten och barnadödligheten i kosovo den högsta i europa - men vi har också en allmän uppfattning om den humanitära katastrofsituationen i kosovo . anser ni inte , herr kommissionär , att detta redan i sig allvarligt skadar vår trovärdighet och tilltron till vår förmåga att leva upp till våra löften ?
och vidare , herr kommissionär , svarar den s.k. humanitära militära insatsstyrkan mot behoven i det katastrofdrabbade kosovo ?
anser ni att man kan rättfärdiga en så stor passivitet , när själva rätten till liv hotas på den europeiska kontinenten ?
jag tror inte att vårt återuppbyggnadsorgan eller insatsstyrkan innan den , vilken har arbetat otroligt hårt i kosovo , skulle anse det vara en riktig beskrivning av deras arbetsinsatser att antyda att de stått bredvid sysslolösa .
jag är säker på att ärade ledamoten inte menade det .
naturligtvis har hon helt rätt när hon säger att unionens trovärdighet står på spel med det som händer inte bara i kosovo utan på hela balkan .
jag är mycket angelägen om att den hjälp vi tillhandahåller anländer snabbt och på ett sätt som ytterligare ökar våra hjälpinsatser .
jag vill endast ta upp två punkter om situationen i kosovo som vi håller på att försöka lösa så positivt som vi kan i överensstämmelse med who .
för det första är jag säker på att ärade ledamoten känner till att under 1990-talet underfinansierade regeringen i belgrad hälsovårdssystemet i kosovo och många albaner upptäckte att de inte fick någon hälsovård alls .
till följd av detta inrättades ett parallellt hälsovårdssystem genom moder teresa organisationen .
vad det således handlar om är inte bara följderna av konflikt utan resultaten av år av misskötsel och ständigt för litet investeringar .
vidare , och jag är säker på att den ärade ledamoten känner till detta likaså , har några av de tragiska historier som man hört från kosovo under de senaste veckorna inte handlat om barndödlighet under graviditet utan barndödlighet efter det att ett friskt barn fötts .
detta gällde fall där kvinnor före eller under fientligheterna tragiskt dödade sina egna barn .
vi har att göra med en fasansfull historia i kosovo .
vi måste arbeta så bra vi kan på hälsovårdsområdet och andra områden för att återställa något som liknar civila normer och civilt uppträdande , men det kommer inte att bli lätt .
herr kommissionär ! jag tackar er för ert svar på den första frågan från min kollega och även på den kompletterande frågan .
jag har dock en del kontakter i kosova och där säger man att de matpaket som delas ut bland annat av echo ofta är av undermålig kvalitet .
i vissa fall har man också hittat insekter och så i maten .
känner ni till det ?
är ni beredd att göra något åt det ?
det är min första kompletterande fråga .
min andra fråga gäller er hänvisning till återuppbyggnaden av sjukhuset i mitrovica .
ni känner kanske till att det sjukhuset ligger i den norra delen av staden och att , med tanke på det spända läget , kosovoalbanerna inte alls får komma in där .
vad gör kommissionen för att se till att även kosovoalbaner får tillgång till sjukhus ?
som svar på den första frågan kommer jag själv att resa till kosovo i början av nästa månad för ett andra besök och jag skall naturligtvis undersöka anklagelsen från ärade ledamoten om echo : s matpaket .
jag har inte hört detta antydas förut , men det är en viktig punkt och jag skall naturligtvis undersöka den när jag är där .
vidare förstår jag inte exakt vad ärade ledamoten menar om mitrovica .
jag var i mitrovica för några månader sedan och såg själv situationen där .
jag förde diskussioner med kommunala ledare från båda sidor , däribland ledaren för den albanska sidan som själv tidigare varit doktor och som var allmänt erkänd för det läkarjobb han hade utfört under fientligheterna och senare .
så jag känner till de mycket allvarliga problem som finns på det sjukhuset och jag kan försäkra den ärade ledamoten att vi kommer att göra allt vi kan för att tillräckliga hälsovårdsinrättningar finns för alla i kosovo , oavsett etnisk grupptillhörighet .
de speciella svårigheterna i mitrovica , exempelvis albanska patienter som har problem att få komma till sjukhus , albansk personal har svårt att få arbeta där - är särskilt akuta problem .
vi skall försöka lösa dem men det är inte lätt .
fråga nr 37 från ( h-0029 / 00 ) :
angående : turkiets blockad mot armenien genom avtalet om partnerskap och samarbete , som undertecknades den 12 oktober 1999 , främjar europeiska unionen aktivt de sociala , ekonomiska och politiska förbindelserna med armenien . vad gör kommissionen för att den turkiska regeringen skall häva den ekonomiska blockaden mot armenien ?
kommissionen stöder varje insats som syftar till att lösa konflikten mellan turkiet och armenien och beklagar att det fortfarande inte har skett någon normalisering av förbindelserna mellan dessa två länder .
under rådande politiska förhållanden är det emellertid orealistiskt att tänka sig att gränsen mellan armenien och turkiet liksom den mellan armenien och azerbajdzjan kan öppnas utan en lösning på konflikten nagorno-karabach .
( de ) herr talman ! kommissionen skall ju också i framtiden föra förhandlingar på grund av anslutningen av turkiet till europeiska unionen .
kommer den att sätta upp som villkor att diskussionen påbörjas först när blockaden här har avbrutits , ty när allt kommer omkring är vi alla grannar , och vi vill ju också vårda grannsämjan inom europeiska unionen ?
jag frågar alltså : kommer kommissionen att göra detta till ett av villkoren för att förbättra de framtida samråden ?
den viktigaste punkten är att stödja insatserna från osse : s grupp i minsk för att hitta en lösning på nagorno-karabach konflikten och vi är beredda att hjälpa till på alla sätt vi kan .
vi har även medverkat på ett omfattande sätt med utvecklingsstöd till armenien inom ramen för tacis-programmet .
låt mitt svar speciellt sättas i samband med frågan om turkiets anslutning till europeiska unionen .
situationen med turkiets förbindelser med dess grannar kommer , såsom den ärade ledamoten begär , att noga granskas inom ramen för strategin för förberedelse för anslutning till unionen .
såsom fastslås i agenda 2000 - och jag citerar : &quot; utvidgning skall inte innebära att gränskonflikter förs in . &quot;
det uttalandet kan inte bli mer tydligt .
men jag upprepar att det viktigaste bidraget vi kan göra är att försöka hjälpa till att lösa den konflikten som har orsakat sådana ekonomiska och humanitära skador .
fråga nr 38 från ( h-0040 / 00 ) :
angående : konsekvenserna av byggandet av ilisudammen i turkiet för de mänskliga rättigheterna med tanke på att turkiet nyligen gavs kandidatlandstatus , vad anser kommissionen om de konsekvenser som byggandet av ilisudammen får för de mänskliga rättigheterna ? detta bygge kommer att medföra en stor omflyttning av den kurdiska befolkningen och av andra invånare i regionen .
kommissionen har ingen information om effekten för befolkningen i regionen av att ilisu- dammen byggs .
vi skall dock överväga att ta upp frågan med de turkiska myndigheterna , tillsammans med andra frågor rörande regional utvecklingspolitik inom ramen för den nya strategin för turkiets förberedelse för anslutning till unionen .
jag har en närbesläktad punkt .
den gäller dammens effekter för tillgång till färskvatten i regionen som helhet .
som ni känner till kommer dammen att begränsa tillgången på vatten till syrien och irak i synnerhet .
med hänsyn till hur ytterst instabil denna region är och många kommentatorers verkligt reella oro över att vi kommer att få se ett ökat antal konflikter , av så kallade &quot; vattenkrig &quot; , under de närmaste decennierna , vad anser kommissionen om den eventuella destabiliserande effekt både i turkiet och i den bredare regionen som denna damm kommer att orsaka ?
kan ni tala om ifall ni verkligen kommer att ta upp även denna fråga ?
vi skall helt klart ta upp den punkt som den ärade ledamoten beskrivit .
vi har fått höra oroliga frågor om detta och jag skall se till att den tas upp .
det har också uttryckts betydande farhågor om den eventuella faran för de arkeologiska lämningarna i området .
vi skall ta upp det också i de framställningar vi gör .
ett antal andra vattenkraftsprojekt som planerats under de senaste 30 åren i turkiet har framkallat oroliga frågor , som följderna för tvångsförflyttade bönder .
på det hela taget verkar dessa ha skötts relativt tillfredsställande och jag hoppas att samma sak kan gälla om detta projekt vilket - för att klargöra frågan - inte är ett projekt i vilket kommissionen deltar i någon form .
vi tackar herr patten för att han har företrätt kommissionen i besvarandet av dessa frågor .
fråga nr 39 från ( h-0036 / 00 ) :
angående : utkastet till en stadga om grundläggande rättigheter det civila samhället ser med tillfredsställelse på utkastet till en stadga om grundläggande rättigheter och förhoppningen är att denna skall kunna anta de utmaningar som europa kommer att ställas inför under det 2l : a århundradet .
kan kommissionen mot denna bakgrund svara på följande frågor :
hur ser kommissionen på innehållet i stadgan ?
vem skall stadgan gälla ?
medborgare i europeiska unionen eller i alla europeiska länder , med tanke på utvidgningen ?
kommer stadgan att befästa europeiska unionens sociala rättigheter eller kommer den att ha en bredare karaktär ?
vilka mekanismer kommer att användas i stadgan för att tydligt säkerställa jämlikhet mellan de båda könen ?
vad anser kommissionen om att införa stadgan i eu-fördraget ?
herr kommissionär ! det är mycket betydelsefullt så här i början av det nya århundradet att europas medborgare , män och kvinnor , uppmanas att ännu en gång definiera sina rättigheter och skyldigheter .
jag hoppas verkligen att detta beslut från rådsmötet i köln skall kunna genomföras .
både globaliseringen och utvidgningen framtvingar en definition av dessa rättigheter .
seattle innebär en verklig källa till problem i detta avseende , och jag hoppas att europeiska rådets möte i nice inte skall innebära ännu ett förlorat tillfälle .
för att medborgarna skall bli delaktiga i denna nya planering , skulle jag vilja veta vad de europeiska organen - närmare bestämt europeiska kommissionen - har för förslag till social och ekonomisk modell för europa under det 21 : a århundradet .
jag har hört era allmänna riktlinjer , och jag skulle vilja fråga er vilken plats barnen , som självständiga individer , har i europeiska kommissionens planering för den nya sociala modellen under det 21 : a århundradet .
jag bör säga er mycket tydligt att , enligt min åsikt och såsom ordförande prodi sade i morse , är utarbetandet av stadgan en politiskt mycket betydelsefull uppgift eftersom den visar att unionen placerar medborgarnas grundläggande rättigheter längst fram bland de politiska angelägenheterna för vårt gemensamma projekts framtid .
inom den ramen måste man klart och tydligt säga på vilka kriterier man grundar sig för att välja rättigheter .
jag tror att det väsentliga kriteriet är medborgarnas rättigheter gentemot de europeiska institutionerna . det är medborgarnas rättigheter såsom de anges i det europeiska projektet som fastställs i unionens fördrag .
jag förstår er omsorg om barnens rättigheter .
jag tror att flera delar av vårt arbete och framför allt av mitt arbete i egenskap av ansvarig för sektorn för rättsliga och inrikes frågor består i att se till barnens rättigheter .
här kommer vi in på ett område där subsidiaritetsprincipen tillämpas fullt ut .
varje medlemsstat har huvudansvaret för att fastställa sitt ansvar gentemot barnen .
när det gäller unionens ansvar som sådant tror jag att barnens rättigheter bör erkännas i stadgan genom att de områden beaktas där unionen kan tillföra ett mervärde till främjandet av den sociala , ekonomiska och till och med , i vidaste mening , medborgerliga situationen för barnen .
jag hoppas att vi kommer att lyckas att anta den utmaning som ledamoten har ställt på kommissionen och på hela konventionen .
herr talman ! jag har haft nöjet att höra kommissionären uttala sig ett antal gånger i denna fråga och jag håller mycket med honom och hans inställning .
jag vill dock ställa en något annorlunda fråga .
vi har just hört kommissionär barnier säga att han är angelägen om att kommunicera bättre med människorna och att inrikta kommissionens informationspolitik mot de större frågor som gemenskapen arbetar med i år .
skulle kommissionären anföra skäl för att någon del av kommissionens informationsbudget används för att informera och samråda med medborgarna i denna fråga om en medborgarstadga ?
det är viktigt att människorna känner sig delaktiga i denna process .
jag vet att själva konventet kommer att bidra mycket på detta område men den har inte de resurser som kommissionen har .
kommer kommissionen att överväga att använda sin informationsbudget för att se till att människor blir intresserade av denna debatt ?
det är kommissionens policy att främja en öppen och bred debatt om stadgan om grundläggande rättigheter , inte bara med icke-statliga organisationer utan också med medborgarna i ett projekt som är så omfattande som stadgan är .
jag kan försäkra er att kommissionen kommer att göra sitt yttersta för att främja debatten om den framtida stadgan om grundläggande rättigheter .
vi kan uppnå det bästa från båda världar genom att få en tydlig text och samtidigt en text som kan användas som ett rättsligt instrument .
det finns ingen motsägelse mellan de två .
vår utmaning är att sammanföra dem i den slutgiltiga versionen av stadgan .
jag är mycket glad att veta att jag kan räkna med ert stöd i denna fråga .
fråga nr 40 från ( h-0095 / 00 ) :
angående : artiklarna 6.1 , 7.1 och 7.2 i fördraget om europeiska unionen i artikel 6.1 i fördraget står det att unionen bygger på principerna om frihet , demokrati och respekt för de mänskliga rättigheterna och de grundläggande friheterna .
av de uttalanden som under de senaste åren gjorts av jörg haider och frihetspartiet framgår det klart att dessa inte respekterar mänskliga rättigheter eller grundläggande friheter för tredjelandsmedborgare och minoritetsgrupper som är bosatta i österrike .
kan kommissionen därför ge besked om när kommissionen tänker åberopa artikel 7.1 om att &quot; en medlemsstat allvarligt och ihållande åsidosätter principer som anges i artikel 6.1 &quot; och yrka på att rådet med kvalificerad majoritet skall fatta beslut om att tillfälligt upphäva vissa av de rättigheter som österrike har till följd av tillämpningen av detta fördrag , inbegripet rösträtten i rådet för företrädaren för österrike ?
herr talman , ärade kollegor ! låt mig börja med att påminna er om kommissionens ståndpunkt när det gäller den nya österrikiska regeringen där ministrar från jörg haiders liberala parti ingår , något som upprepades i morse av ordförande prodi .
jag syftar givetvis på kommissionens uttalande från den 1 februari 2000 och vars huvudpunkter jag vill börja med att påminna om .
kommissionen försäkrade på nytt och försäkrar i dag igen att man delar den underliggande oron i det portugisiska ordförandeskapets uttalande från den 31 januari .
oron är berättigad och skälig .
vi behöver inte påminnas om jörg haiders politiska bana och hans otaliga offentliga uttalanden , främlingsfientliga och rasistiska , med andra ord antieuropeiska .
att ett klart extremistiskt , rasistiskt och främlingsfientligt parti kan komma till makten i en av europeiska unionens medlemsstater är något som de övriga deltagarna i det europeiska projektet inte kan sluta att oroa sig över , på samma sätt som det inte är likgiltigt för europeiska kommissionen .
för det andra så upprepade kommissionen , och upprepar igen , sitt åtagande att fortsätta fullgöra sina skyldigheter som fördragens väktare , särskilt det som åsyftas i artikel 6 och 7 i eu-fördraget .
en av de viktigare reformerna i amsterdamfördraget var just de grundläggande principernas tydlighet , vilket är medlemsländernas gemensamma arv och institution för den kontrollapparat som krävs för att se till att de åtföljs och att en reaktion sker om någon av principerna kränks .
kommissionen visade därmed i praktiken sin tillgivenhet för en av de grundläggande principerna : rättsstatens .
en sådan princip ålägger kommissionen att hålla sig inom de gränser som fastställts genom fördragen och det är i det här sambandet som uttalandet från den 1 februari skall ses .
kommissionen är inte en stat , den varken kan eller bör agera som om den vore det .
men för att besvara ledamotens fråga vill jag påminna om att den mekanism som instiftats i artikel 7.1 i eu-fördraget för att aktiveras kräver en bekräftelse på , jag citerar , &quot; att en medlemsstat allvarligt och ihållande åsidosätter principer i artikel 6 &quot; .
jag upprepar , ett allvarligt och ihållande åsidosättande är ett oumbärligt villkor för att kommissionen skall kunna uppmana rådet att vidtaga åtgärder mot ett medlemsland .
för mig är det uppenbart att villkoren inte är uppfyllda för att tillämpa dem på situationen i österrike .
jag tror inte att jag misstar mig när jag säger att vi alla hoppas att ett sådant allvarligt och ihållande åsidosättande av de mänskliga rättigheterna och demokratin aldrig någonsin kommer att inträffa , varken i samband med österrike eller något annat land inom unionen .
jag vill dock försäkra er alla här i dag att min personliga ambition och kommissionens , som ordförande prodi bekräftade i morse , är att göra allt som står i vår makt för att det inte skall bli nödvändigt att tillämpa artikel 7 .
jag vill emellertid också säga att vi inte kommer att tveka att använda den om det behövs .
de värden som står på spel är alldeles för viktiga och grundläggande för att visa hänsyn eller kompromissa . §
§ människor och regeringar bör värderas mera efter vad de gör än vad de säger .
i fallet med österrike är uttalandena åtminstone motsägelsefulla .
å ena sidan kan vem som helst av oss samla ihop ett antal upproriska meningar från det österrikiska liberala partiet .
å andra sidan upprepar den nya österrikiska regeringen i sitt program sin ambition att försvara demokratin och de mänskliga rättigheterna .
inom kort får vi ett ypperligt tillfälle att se vilken av de här två sidorna som är den rätta .
jag tänker här på vilken ståndpunkt den österrikiska regeringen kommer att inta i rådet beträffande kommissionens förslag om ett åtgärdsprogram för kampen mot diskriminering samt två direktiv .
ett som tillämpar principen om alla människors rätt till lika bemötande oavsett ras eller etniskt ursprung och ett annat som erbjuder ett skydd mot diskriminering vid anställning på grund av ras eller etniskt ursprung , religion och sexuell inriktning .
det är relevanta dokument som godkänts i enlighet med artikel 13 i fördraget och där gemenskapen ges fullmakt att bekämpa diskriminering grundad på ras , etniskt ursprung , kön osv.
låt mig avslutningsvis försäkra ledamoten om att kommissionen kommer att fortsätta att vara vaksam och vi kommer inte att sluta fullgöra våra skyldigheter , om detta skulle visa sig vara nödvändigt .
jag tackar kommissionären för hans svar på min fråga .
men är kommissionär vitorino medveten om inte bara haiders och frihetspartiets uttalanden utan också deras gärningar ?
haider har i själva verket varit verksam i ledningen i den södra provinsen kärnten där han har lett en rasistisk och främlingsfientlig kampanj mot den slovensktalande minoriteten i den regionen som är österrikiska medborgare , där han har försökt att avskaffa tvåspråksutbildningen och där det har det skett en klar diskriminering mot romerbefolkningen och immigrantbefolkningen .
kan kommissionären besvara två frågor .
för det första talade han om bekräftelse .
kan han tala om hur den bekräftelsen skall ske och vem som skall göra den ?
för det andra , håller han inte med om att ifall den nuvarande regeringen på nationell nivå skulle bedriva den slags politik som haider och frihetspartiet bedrivit på regional nivå det klart skulle strida mot artikel 6.1 i fördraget i fråga om grundläggande fri- och rättigheter och det skulle falla på kommissionen att vidta nödvändiga åtgärder ?
vi talar inte om uttalanden här .
vi talar om gärningar av frihetspartiet och haider .
jag anser det helt klart att det är kommissionens ansvar att noggrant följa utvecklingen av situationen i medlemsstaterna i enlighet med de förfaranden och normer som inryms i artikel 6 och som berättigar tillämpning av artikel 7 i fördraget .
därför är jag helt förvissad om att kommissionen mycket noga kommer att kunna följa utvecklingen av situation i österrike liksom i många andra medlemsstater .
om något konkret fall av ständig kränkning av de mänskliga rättigheterna begåtts av regeringen i en medlemsstat kommer vi att var helt i stånd att reagera och agera därefter .
jag förlitar mig inte bara på samarbetet från europaparlamentets ledamöter utan även på samarbetet från icke-statliga organisationer som alltid har lämnat ett viktigt bidrag till kommissionens politik mot diskriminering .
beträffande situationen i kärnten , måste vi undersöka den närmare .
ärade ledamoten tog upp frågan .
skyddet för etniska minoriteter och för minoriteter som talar en särskilt språk är ett del av programmet och i de två direktiv som kommissionen har lagt fram för rådet .
vi bör inte enbart inrikta denna debatt på den österrikiska frågan .
den frågan kräver eftertanke , debatt och om så krävs , åtgärd .
jag hoppas uppriktigt att alla medlemsstater skall ta möjligheten i fråga om denna handlingsplan och dessa två direktiv som kommissionen lagt fram för rådet att upprepa i klara och konkreta termer deras godkännande av handlingsplanen och direktiven och deras åtagande att bekämpa diskriminering , rasism och främlingsfientlighet varhelst det kan tänkas ske .
tack så mycket , herr vitorino , för ert värdefulla bidrag till frågestunden .
frågor till wallström
fråga nr 41 från ( h-0021 / 00 ) :
angående : elektriskt och elektroniskt avfall för varje år som går står eu inför en allt större mängd elektriskt och elektroniskt avfall ( 6 miljoner ton 1998 ) som framför allt beror på apparaterna blivit föråldrade i allt snabbare takt .
miljöproblemen till följd av att dessa apparater förbränns eller slängs på soptippen beror i främsta rummet på att de innehåller farliga ämnen ( bly , kadmium , kvicksilver , hexavalent krom , pvc och halogenerade flamskyddsmedel ) .
ett utkast till förslag till direktiv i syfte att reglera administrationen av dessa avfall gav upphov till tre på varandra följande versioner , den senaste från juli 1999 .
kan kommissionen förklara varför administrationen av det här projektet tagit så tid , trots att det i princip borde ha varit klart 1998 ?
stämmer det att den amerikanska regeringen motsätter sig de flesta bestämmelser i det nuvarande förslaget och att den till och med hotar att dra eu inför wto ( för brott mot artikel xi i gatt-avtalet och artikel 2.2 i avtalet om tekniska handelshinder ) ifall förslaget antas ?
kommissionen håller med parlamentsledamoten om att den nuvarande hanteringen av elektriskt och elektroniskt avfall inom europeiska unionen orsakar betydande miljöproblem .
kommissionen har därför beslutat att utarbeta ett förslag i ämnet och har sedan 1997 tagit upp frågan med alla berörda parter .
resultaten från denna debatt och de grundliga efterforskningar som görs på området granskas nu av kommissionen .
vissa delar av förslaget har utsatts för kritik , bland annat utfasningen av vissa tungmetaller och bromerade flamskyddsmedel samt tillämpningen av principen om tillverkarens ansvar för hanteringen av elektriskt och elektroniskt avfall .
förenta staternas delegation vid europeiska unionen har ställt sig tveksam till några punkter i det senaste samrådsdokumentet , bland annat just utfasningen av ovannämnda ämnen och vissa frågor som gäller principen om tillverkarens ansvar .
förenta staternas huvudargument i detta sammanhang är att de ifrågavarande bestämmelserna påstås vara oförenliga med internationell handelsrätt .
kommissionen har för närvarande delegationens argument under övervägande .
låt mig tillägga att mina planer är att före påsk för kommissionen kunna presentera ett förslag om hantering av elektriskt och elektroniskt avfall .
min fråga gällde just den amerikanska regeringens reaktion på texten i det förberedande projektet .
det finns nämligen tre förberedande texter och den sista enligt min vetskap från juli 1999 .
är det således denna text som ni skall lägga fram eller en ändring i förhållande till den ursprungliga versionen ? .
den tredje versionen var nämligen redan svagare än den andra versionen till följd av den amerikanska industrins anmärkningar , som följdes upp av den amerikanska regeringen .
jag vill i synnerhet påpeka att , när ni talar om den internationella rätt med vilken det sägs att texten inte överensstämmer , syftar ni nämligen på världshandelsorganisationens regler .
den amerikanska regeringens påståenden gäller det faktum att det skulle vara att gå emot wto : s regler att på sikt förbjuda förekomsten av farliga ämnen i elektriskt och elektroniskt avfall .
det bekymrar mig personligen eftersom det skulle betyda att om man antar en text står man ständigt under hot om en attack inför världshandelsorganisationen , och det försvagar således fullständigt den europeiska miljölagstiftningen , i synnerhet detta förslag .
tack för följdfrågan .
det är viktigt att jag får tillfälle att svara på den .
det är klart att i en process som denna , där vi diskuterar en mycket stor avfallsström i europa av både elektriskt och elektroniskt avfall , pågår en ständig dialog mellan olika inblandade parter .
vi har haft en bra dialog och har utvecklat ett förslag under processens gång .
vissa avsnitt har stärkts , andra har vi kanske fått kompromissa litet för mycket med .
vi håller fortfarande på att skriva på texterna , och dialogen med de olika inblandade parterna pågår ända in i sista minuten .
jag vill säga att jag inte anser att förenta staternas inblandning i denna fråga skall låta oss styras på ett sådant sätt att vi inte tar tillräcklig miljöhänsyn .
jag värjer mig verkligen mot att man ständigt skall kunna hänvisa till wto och handelsregler för att förhindra att vi i eu skaffar oss radikala miljöbestämmelser .
min utgångspunkt är att vi skall göra det .
jag är emellertid beredd att lyssna på alla argument .
jag har exempelvis nyligen träffat företrädare för elektronikbranschen . de lämnade förslag - också praktiska - till hur man skulle kunna förbättra vårt förslag .
jag vill dock bestämt tillbakavisa påståendet att jag skulle låta förenta staterna styra utformningen av vårt direktiv .
det är faktiskt så att jag menar att vi måste visa vägen , vilket också kommer att prägla det slutgiltiga förslaget .
fråga nr 42 från ( h-0026 / 00 ) :
angående : gender och miljö så gott som samtliga aktörer i rio- och kyotoprocesserna - enskilda organisationer , medborgarrörelser , regeringar världsbanken , fn och hjälporganisationer - ansåg att kvinnor i högre grad skall delta i beslutsfattande inom miljöområdet.fler kvinnor i beslutsfattande positioner inom olika miljöorgan gör att de förhärskande manliga referensramarna utvidgas till att omfatta inte bara frågor som berör företagande utan även sociala rättvisefrågor .
är kommissionen beredd att anta en handlingsplan för att öka kvinnors aktiva deltagande i beslutsfattande även inom miljöområdet .
kommissionen har sedan 1988 ett handlingsprogram för lika möjligheter för kvinnor och män .
med hjälp av det nuvarande programmet , som omfattar åren 1997 till 2000 , försöker man utveckla en arbetskultur , som innebär att både manliga och kvinnliga värden integreras , och att hänsyn tas till könsspecifika behov .
ett av programmets syften är att utarbeta och övervaka metoder , strategier och åtgärder , som främjar en jämn könsfördelning i beslutsprocessen , däribland på högre befattningar .
inom ramen för detta handlingsprogram utarbetar varje enskilt generaldirektorat en särskild åtgärdsplan .
ett av målen i åtgärdsplanen är att öka antalet kvinnor i ledande ställning .
den nya kommissionen har som mål att fördubbla antalet kvinnliga chefer under sin mandatperiod .
denna linje drivs särskilt aktivt på generaldirektoratet för miljö , där för närvarande 60 procent av direktörerna och 20 procent av enhetscheferna är kvinnor .
vår politik är att gynna rekryteringen av kvinnor till administrativa tjänster för att skapa en reserv av lämpliga kandidater för framtida chefstjänster .
för närvarande är 24,5 procent av våra a-tjänstemän kvinnor . vi hoppas att antalet kommer att öka stadigt .
vi anstränger oss dessutom för att locka kvalificerade kvinnor att delta i de samrådsforum som vi organiserar .
när det gäller våra externa partners kan vi bara föregå med gott exempel och uppmuntra deras ansträngningar att demokratisera sina beslutsprocesser .
när det gäller mer allmänna frågor om integrering av jämställdhetsperspektivet , känner ni säkert till att denna princip ingår i amsterdamfördraget .
i artikel 3 i fördraget anges att gemenskapen i all verksamhet som avses i denna artikel skall syfta till att undanröja bristande jämställdhet mellan kvinnor och män och att främja jämställdhet mellan dem .
kommissionen ger sitt fulla stöd till ansträngningarna på detta område och håller på att undersöka om specifika åtgärder kan vidtas på miljöområdet .
naturligtvis vill jag passa på att säga att jag uppskattar den roll som europaparlamentets kvinnoutskott , och inte minst dess ordförande , spelar .
låt mig bara påminna om att när den nuvarande kommissionen så småningom godkändes fick varje kommissionär en fråga från kvinnoutskottet om hur de inom just sitt verksamhetsområde skulle sköta jämställdheten .
vi kommer noggrant att granska varje kommissionär , så jag vill härmed förvarna även de andra kommissionärerna .
tack så mycket för svaret !
jag tolkar det faktiskt som ett ja till att det är en handlingsplan som behövs - en handlingsplan för att få fler kvinnor att delta inom specifika miljöområden .
låt mig också säga att pekingdeklarationen understryker vikten av att ha institutionell kapacitet för att ta med ett jämställdhetsperspektiv i all miljöprogrammering .
miljöinstitutioner saknar ofta kunskaper och procedurer för att inkorporera ett sådant perspektiv i sitt dagliga arbete .
jag vill naturligtvis veta om kommissionären är villig att integrera jämställdhetstänkandet i miljöpolitiken och i miljöprogrammen .
om hela politiken skall genomsyras , tror jag att det är särskilt viktigt att cheferna på hög nivå har denna grundläggande kunskap .
naturligtvis är min bild av mainstreaming att detta måste prägla allt vi gör .
i den plan som utarbetas på mitt generaldirektorat spelar jämställdhetsfrågorna en mycket viktig roll .
jag är också beredd att själv gå in och exempelvis leda seminarier i ledarskap eller andra ämnen för att uppmuntra kvinnor att ta på sig vidare uppgifter inom kommissionen .
om vi skall kunna motivera alla , tror jag att det är väldigt viktigt att detta budskap sänds hela vägen uppifrån och ned - eller nedifrån och upp om du så vill .
min bild av miljöarbete i stort är att det många gånger domineras av kvinnor .
det handlar om att detta måste fortplantas , så att kvinnor har en chans att också få chefsjobb eller komma till högre positioner inom miljöarbetet .
jag vill påstå att vår åtgärdsplan avspeglar detta , men den kan säkert göras bättre .
jag har en viss erfarenhet av att upprätta planer och följa upp dem .
jag hoppas att detta skall komma till nytta .
fråga nr 43 från ( h-0045 / 00 ) :
angående : området vid mynningen av floden boyne och företaget drogheda området vid mynningen av floden boyne är klassificerat som ett särskilt skyddsområde enligt direktivet om vilda fåglar och man överväger för närvarande att klassificera det som ett särskilt bevarandeområde enligt habitatdirektivet på grund av dess internationella betydelse .
marindepartementet , grevskapsrådet i louth och företaget drogheda har godkänt uppförandet av en ny hamn i det särskilda skyddsområdet och till och med avskaffandet av en strandremsa i stegrennan , som nyligen införlivades i det särskilda skyddsområdet på kommissionens uttryckliga uppmaning .
dessutom har man uppfört ett mycket stort lagerhus . det har visat sig vara svårt att få tag på byggnadstillståndet för detta lager , och drogheda planerar samtidigt annan infrastruktur .
hur kan kommissionen säkerställa att sådana projekt som finansieras via strukturfonderna inte går stick i stäv mot miljöskyddsbehoven i området ?
är kommissionen beredd att inställa finansieringen helt och hållet i väntan på att utvecklingsplanerna för detta område skall ses över ?
kommissionen känner till uppförandet av hamnen , men vet inget om det lagerhus , eller den övriga infrastruktur som parlamentsledamoten nämner .
hamnens uppförande får stöd från strukturfonderna och medför i huvudsak att utloppet i floden boynes mynning muddras och att muddermassorna mellanlagras på stegrennans strandremsa .
floden boynes mynningsområde är klassificerat som särskilt skyddsområde enligt direktivet om vilda fåglar .
detta innebär att man vid all exploatering i eller vid boynesmynningen , som kan komma att påverka det särskilda skyddsområdet , måste beakta de skyddsbestämmelser för området som fastställts i gemenskapens habitatdirektiv .
sedan 1998 har det till kommissionen kommit in ett antal klagomål , där man hävdar att hamnanläggningen kommer att skada stegrennans strandremsa , som numera ingår i det särskilda skyddsområdet , och att man inte har beaktat de relevanta skyddsbestämmelserna .
efter att ha granskat dessa klagomål under 1998 och i början av förra året - projektet erhöll under denna tiden inga medel från strukturfonderna- blev kommissionen på sommaren 1999 övertygad om att man vid uppförandet av hamnen hade beaktat de relevanta skyddsbestämmelserna .
en detaljerad miljökonsekvensbedömning hade gjorts .
den mest negativa följden av projektet , förlusten av stegrennans strandremsa , skall endast vara tillfällig , och entreprenören är skyldig att helt återställa strandremsan .
på kommissionens uppmaning införlivades stegrennansstrandremsa formellt i boynesmynningens särskilda skyddsområde , från vilken den tidigare hade varit utesluten .
för att uppväga de negativa effekterna av strandremsans tillfälliga försvinnande på berörda fågelpopulationer var det dessutom meningen att andra livsmiljöer i mynningsområdet skulle förbättras .
sedan sommaren förra året har emellertid den sistnämnda åtgärden varit omtvistad .
först drog de irländska myndigheterna tillbaka sitt tidigare förbättringsåtagande .
de förnyade sedan sitt åtagande efter det att en icke-statligt irländsk miljöorganisation hade anfört klagomål inför irländsk domstol .
det nya åtagandet innehöll dock smärre ändringar , som i sin tur ledde till ytterligare ett klagomål .
mot bakgrund av att irland har åtagit sig att vidta kompensationsåtgärder , och med tanke på att andra frågor redan har lösts , vill kommissionen för närvarande inte föreslå att man ställer in finansieringen från strukturfonderna .
kommissionen vill dock reda ut spörsmålet om kompensationsåtgärden avseende förbättrade livsmiljöer med de irländska myndigheterna , särskilt i ljuset av den ännu oavslutade processen inför irländsk domstol .
jag förstår inte riktigt det som kommissionären sade .
den gyttjiga strandremsan vid stregrennan , som gjordes till ett särskilt skyddsområde på kommissionens begäran har förstörts helt i detta skede .
det är uppenbart att de aktiviteter som har skett där klart bryter mot eg-direktiven .
ni säger att det inte kommer att anslås mer medel .
jag skulle vilja veta om ni tänker stoppa finansieringen helt i detta skede tills det blir en ordentlig utredning .
om inte , varför inte ?
om ni tänker göra det , när exakt kommer ni att göra det ?
är det rätt och lämpligt att det departement som äger företaget också är den myndighet som utfärdar tillståndet och även den myndighet som praktiskt taget tar emot pengarna från eu och ger det till ett företag som det äger till 100 procent ?
är detta rätt och lämpligt ?
vad anser ni om det ?
varje bidrag från eu till projektet måste stoppas eftersom det klart bryter mot eg-direktiven .
även det område som utsetts som särskilt skyddsområde av kommissionärerna har förstörts .
skadestånd efteråt kan inte gottgöra den skada som uppstått .
den första rättsliga utmaningen kom efter det att arbetet med att uppföra hamnen inletts tidigt på hösten 1999 utan att förbättringar i form av kompenserande livsmiljöer inrättats .
till följd av det gick de irländska myndigheterna med på att på nytt börja avlägsna marskgräset men denna gång på mekanisk väg .
användningen av mekaniska hjälpmedel ledde till ytterligare ett klagomål - det är vad jag tog upp även i mitt första svar - grundat på argumentet att man genom mekaniskt avlägsnande skulle skada underliggande gyttjemark och orsaka ekologiskt skadlig spridning av marskgräset i flodmynningen .
det finns hittills inget slutgiltigt resultat på detta klagomål .
beslut om nödvändiga kompensationsåtgärderna är en fråga för de nationella myndigheterna och kräver inget föregående godkännande av kommissionen .
kommissionens roll är att se till att de normer som gäller enligt fågeldirektivet beaktas fullt ut och uppenbarligen skulle det bli problem med kompensationsåtgärder som i sig själva orsakar skada .
i detta fall föreslår kommissionen att få ytterligare klargöranden från de irländska myndigheterna om det aktuella läget med kompensationsåtgärderna och eventuella problem med det mekaniska avlägsnandet av marskgräs .
vi är för närvarande inte beredda att föreslå att man ställer in finansieringen från strukturfonderna .
herr talman ! tyvärr är det speciella fall som mckenna tog upp inte ett isolerat sådant .
det finns andra exempel på naturskydd på särskilda vetenskapliga områden där skador uppstått till följd av finansiering från eu .
kommer kommissionen att överväga att utfärda föreskrifter till alla medlemsstater om att om den i framtiden upptäcker att man bryter mot de europeiska miljödirektiven eller tillämplig miljökonsekvensbedömning inte skett kommer den inte bara att inställa vidare finansiering utan även att upphäva beslut om redan beviljade medel , med andra ord , återkräva pengar från medlemsstaterna ?
det är endast en sådan åtgärd som kommer att avskräcka denna praxis i framtiden .
som europaparlamentarikerna säkert känner till , gick det under förra året ut ett gemensamt brev från våra föregångare i kommissionen , ritt bjerregaard och monika wulf-mathies angående förhållandet mellan strukturfonderna , pengar från strukturfonderna och skyddet i habitat- och fågeldirektiven .
det budskap som sändes ut i detta gemensamma brev gäller fortfarande .
vi kan inte med ena handen dela ut pengar och med den andra dra länderna inför domstol och kanske så småningom få böter utdömda .
det är därför viktigt att detta står i samklang .
naturligtvis kan svåra avvägningsfall bli följden .
som jag ser det , är dock den främsta effekten att länderna tänker sig noga för och framför allt ser till att skicka in sina listor över natura 2000-platser , så att vi har möjlighet att övervaka och följa upp på ett ordentligt sätt .
där brister irland i likhet med andra medlemsländer , men vi hoppas att vi skall kunna se resultat av denna påtryckning .
jag vill ännu en gång påpeka att det som stod i detta brev fortfarande är giltigt .
det tillåter inte arbetsordningen .
ni får lov att diskutera det utanför plenisalen , fru ledamot .
frågor till barnier
fråga nr 44 från ( h-0020 / 00 ) :
angående : partnerskap och den tredje gemenskapsstödramen i grekland den nya förordningen ( eg ) 1260 / 1999om allmänna bestämmelser för strukturfonderna betonas , i motsats till i föregående förordning , att partnerskap skall förstärkas och att regionala , lokala och övriga behöriga offentliga myndigheter , arbetsmarknadens parter , näringslivets organisationer och alla andra relevanta organ skall delta i att förbereda och finansiera , övervaka och utvärdera stödåtgärder .
enligt upprepade klagomål från lokala myndigheter är förfarandena vad gäller den nya grekiska gemenskapsstödramen dock oförändrade och &quot; parternas &quot; roll framhävs inte alls . kan kommissionen , mot denna bakgrund , svara på följande frågor :
har den grekiska regeringen tillfogat några ändringar till förfarandena för att bredda partnerskapens sammansättning så att dessa i synnerhet även omfattar lokala myndigheter och andra representativa organ ?
vad innebär vidare de lokala myndigheternas ökade roll i förberedelsen och finansieringen av den tredje gemenskapsstödramen ? vilka åtgärder kommer slutligen kommissionen att vidta för att säkerställa ökat deltagande från &quot; parternas &quot; sida inom alla förfaranden som den nya gemenskapsstödramen omfattar ?
tillåter ni mig att förlänga margot wallströms svar till ordförande david martin med en mening för att säga att eftersom det handlade om en gemensam skrivelse mellan våra båda föregångare anser jag i egenskap av efterträdare till wulf-mathies att skrivelsen förvisso fortfarande är giltig och att jag i gott samförstånd skall ta itu med att tillsammans med margot wallström kontrollera om de projekt som finansieras genom strukturfonderna är förenliga med eu : s miljödirektiv och -politik .
det är också en före detta miljöminister som svarar er , ordförande martin .
jag skulle nu bara vilja säga några ord till alavanos som förlåter mig denna inträngning i ett annat ämne för att säga till svar på hans fråga att kommissionen inom ramen för förberedelsen av den nya programplaneringsperioden förvisso har sett till och kommer att se till att partnerskapsprincipen tillämpas .
jag tillåter mig att här påminna om , men ni vet det , att anslutningen av de regionala och lokala myndigheterna till gemenskapens verksamhet utgör en av de främsta beståndsdelarna i den nya förordningen för strukturfonderna från berlin .
när det mer speciellt rör tillämpningen av partnerskapsprincipen vad gäller den kommande gemenskapsstödramen i grekland har kommissionen kunnat notera att de offentliga myndigheterna i stor utsträckning har fått bidra till utarbetandet av den grekiska planen för regional utveckling för perioden 2000-2006 .
alavanos vet att jag för övrigt har varit där två gånger under ganska tragiska omständigheter till följd av jordbävningsdramat och under dessa besök har jag kunnat diskutera med den grekiska regeringen och påminna om angelägenheten att beakta partnerskapsmålet och -kravet .
när det gäller följande faser , herr ledamot , det vill säga utarbetandet av de nationella och regionala programmen räcker det inte att detta mål beaktas på nationell och teoretisk nivå , det måste göras konkret i de program som utgår från gemenskapsstödramen på de nationella , regionala och lokala planen .
när det gäller uppföljning och förvaltning av programmen har jag ännu inte i detta ögonblick mottagit de nationella bestämmelser som föreslagits av den grekiska regeringen för tillämpning av artikel 8 i den nya förordningen .
jag kan meddela er att jag , inom ramen för förhandlingarna om den tredje gemenskapsstödramen som för närvarande pågår , har bett att bestämmelserna i samband med partnerskapsprincipen skall respekteras fullt ut , inbegripet för de regionala och lokala myndigheterna och inbegripet för allt som rör icke-statliga organisationer och sammanslutningar .
denna princip bör sålunda överföras inom ramen för den tredje gemenskapsstödramen , i synnerhet genom deltagande av samtliga partner till uppföljningskommittén .
herr ledamot , det är det svar jag kan ge er .
jag tackar kommissionären . jag ifrågasätter inte alls hans avsikter och insatser som rört sig i en positiv riktning .
men situationen är helt annorlunda .
just nu får vi uppleva en stark maktkoncentration och både statlig och partipolitisk maktberusning när det gäller bidragen från europeiska unionen .
jag kan inte förmedla tv-programmen här , men jag har tagit med mig några grekiska tidningar till er från veckorna före valet .
i alla greklands söndagstidningar kan man läsa : ministeriet för offentliga anläggningsarbeten om strukturfonden : tack vare ministern ; jordbruksministeriet : tack vare jordbruksministern - några veckor före valet - telekommunikationsministeriet : tack vare telekommunikationsministern ; utbildningsministeriet : tack vare utbildningsministern och så ett fotografi på ministern ; arbetsmarknadsministeriet : tack vare arbetsmarknadsministern , ett fotografi på ministern och ett på biträdande ministern och bakom allt detta emblemet för gemenskapens strukturfonder .
vi har bara några veckor kvar till valet .
propaganda för parti och kandidater , som finansieras med hjälp av gemenskapens strukturfonder .
jag ställer en fråga till kommissionären : kommer kommissionen att tiga ?
kommer kommissionen att ta upp det här med den grekiska regeringen , eller kommer denna kommission att utvecklas i samma patologiska riktning som den föregående ?
herr alavanos , jag har förstått att ni kastar de dokument åt vänster som ni har nämnt .
det skulle vara mig ett nöje om vi ville ge mig dem så att jag kan läsa dem - ja , jag kommer att låta översätta dem - och att jag tittar på vad som liknar information , kommunikation , som jag bara kan glädja mig åt i egenskap av kommissionär med ansvar för regionalpolitik , och propaganda .
och därefter om det är absolut nödvändigt att jag gör det kommer jag att lämna synpunkter eller rekommendationer till den grekiska regeringen .
jag skulle således bli mycket lycklig , herr ledamot om ni kunde ge mig dokumenten eller också går jag och hämtar dem om en stund på golvet i er grupps rad .
därmed sagt att jag trodde att er fråga mer avsåg partnerskapet .
bortom dessa frågor förbundna med den förberedande valperioden som ni anger , säger jag än en gång att jag är bekymrad över att de regionala och lokala myndigheterna är anslutna på samma gång som icke-statliga organisationer .
men jag kan inte heller skriva något annat än det som står i den allmänna förordningen om strukturfonderna och anger att kommissionen skall arbeta med medlemsstaternas regeringar och att det är den grekiska regeringen som jag har till partner , såsom första partner .
sedan måste jag försäkra mig om att partnerskapet sprids , eftersom jag är decentraliserad skall jag försäkra mig om det .
jag kan inte göra annat än att arbeta med den grekiska regeringen .
jag tror att vår kollega alavanos kommer att ge kommissionsledamoten alla dessa uppgifter , så att han kan ta ställning till dem , för det är faktiskt fråga om propaganda och inte något slags reklam för gemenskapens program .
men i själva sakfrågan vill jag be kommissionären att ta hänsyn till följande : att grekland i fråga om samtliga både nationella och regionala program betraktas som en enda region som - i partnerrelationen till europeiska unionen ­ företräds av centralförvaltningen , av centralregeringen .
detta innebär att varken de lokala självstyrelseorganen eller - än mindre - icke-statliga organisationer , som t.ex. de jordbrukskooperativa företag som skulle kunna vara intresserade av en utveckling av jordbrukssektorn , deltar i utarbetandet av förslag i fråga om gemenskapens tredje stödprogram och inte heller har medverkat i fråga om gemenskapens tidigare stödprogram .
hur kan kommissionen hantera denna fråga ?
än en gång theonas , säger jag om vad jag sade till alavanos , jag kommer att nära titta på och , om det behövs , kommer jag att inom ramen för och med iakttagande av strukturfondernas förordning lämna synpunkter på den användning man gör , inte av strukturfonderna som ännu inte har använts utan om förhandlingen före tilldelningen av dessa strukturfonder .
men än en gång , jag måste respektera den nationella myndighet med vilken jag skall genomföra förhandlingen .
jag kommer ändå att se det hela på ett objektivt sätt .
herr theonas , om ni har rekommendationer eller förslag om anslutning av den ena eller andra strukturen - ni talade om kooperativ om jag förstod rätt - är jag öppen och jag är beredd , på grundval av förslag från europaparlamentets ledamöter , ni har er roll och jag har min , att ta över förslag så länge de respekterar tanke och innehåll i förordningen om strukturfonderna .
varför skulle jag inte säga att vi från den grekiska regeringens sida tidigare år har noterat vissa brister när det gäller tillämpningen av den nya förordningen och den föregående förordningen om anslutning av företrädare för det civila samhället .
jag säger det objektivt och när man upptäcker ett problem eller brister måste man avlägsna problemet eller bristerna .
jag skall således se till att det blir gjort inom ramen för genomförandet av den nya gemenskapsstödramen .
fråga nr 45 från ( h-0041 / 00 ) :
angående : finansiering från strukturfonderna av forskning på kärnkraftsområdet kan kommissionen bekräfta att det i den senaste programperioden för strukturfonderna , 1994-1999 , inte utgick något stöd till forskning inom kärnfusion och kärnfission ?
kan den också vid de pågående förhandlingarna med medlemsstaterna om planer och program för den nya perioden , 2000-2006 , arbeta för att inte bevilja några finansieringsåtgärder för den här typen av forskning ?
vilken roll kommer å andra sidan strukturfondsstödet att spela för att främja förnybara energikällor ?
kan man förvänta sig att finansieringen från strukturfonderna inom energipolitiken inriktas på att främja regionala och förnybara energikällor ?
kommer stöd från strukturfonderna även att utgå till de stora näten för energiöverföring ? ¿
jag skulle vilja svara isler béguin på den första punkten och påminna henne om att förbättringen av den vetenskapliga grunden och regionernas tekniska kapacitet i syfte att öka konkurrensförmågan utgjorde en av gemenskapens prioriteringar under den föregående programplaneringsperioden .
det stöd som tilldelas genom strukturfonderna till förmån för teknisk sammanhållning , det vill säga forskning och teknisk utveckling vad gäller gemenskapsstödramarna under denna period uppskattas till omkring 7,5 miljarder euro .
det är ungefär 6 procent av det sammanlagda gemenskapsbidraget , fru ledamot .
vad beträffar just ert bekymmer vill jag säga er att liksom under den föregående perioden har kommissionen inte för avsikt att direktfinansiera forskning och teknisk utveckling på området för fusion eller fission i samband med kärnkraft genom strukturfonderna .
det fortsätter att vara på medlemsstaternas förvaltningsmyndigheters ansvar att välja de projekt som genomförs inom ramen för dessa gemenskapsstödramar .
fru ledamot , även om det inte utgör en prioritering för gemenskapen kan en medlemsstat besluta att finansiera projekt för forskning och utveckling på den civila kärnkraftens område så länge som dessa projekt bidrar till den regionala utvecklingen och utan att för den skull systematiskt informera kommissionen om det .
när det gäller er andra punkt , som ni vet intresserar mig och fortsätter att intressera mig i hög grad , de förnybara energierna , läggs kommissionens tillnärmning fram i dokumentet om strukturfonderna och deras samordning med sammanhållningsfonden .
de avser att investeringar inom sektorn för förnybara energier bör uppmuntras eftersom de främjar utveckling av lokala resurser där de bidrar till beroendeminskning i förhållande till energiimport och är också sysselsättningsskapande på lokal nivå .
jag har kunnat kontrollera det , till exempel vid ett besök i portugal för några dagar sedan på azorerna , där det handlar om en naturlig källa till förnybar energi .
strukturfondernas bidrag till förmån för en större genomträngning på marknaderna av förnybara energier , underströks också i kampanjen för säljstart för förnybara energikällor som inletts av generaldirektoratet för transport och energi .
när det slutligen gäller de stora energinäten , avses också i riktlinjerna ett finansiellt deltagande genom fonden för utveckling av transportnät för energi , när denna bidrar till att minska beroendet gentemot en extern leverantör eller för att bekämpa isoleringseffekter .
det gäller i synnerhet för den region som jag nämnde , azorerna , men också för samtliga områden i de yttersta randområdena och , jag vill tillägga , också för vissa regioner som är handikappade genom isolering på grund av berg , till exempel .
jag har hört ert svar men , å andra sidan , om jag ställde frågan är det just för att vi är oroliga , eftersom ett projekt kallat &quot; international thermonuclear experimental reactor &quot; förekommer inom ramen för betänkandet om den tredje gemenskapsstödramen för forskning .
det uppgår till flera miljarder euro och områden som kan få strukturfonder , såsom mål 1-områdena , skulle kunna få ta emot denna typ av anläggning .
det som vi skulle vilja veta , det är nämligen om kommissionen skulle vara beredd att finansiera denna typ av projekt inom ramen för anläggningen av denna forskningsplats och kanske inte direkt inom den specifika ramen för &quot; kärnforskning &quot; .
herr barnier , förlåt mig men ni svarade inte helt och hållet på den andra delen av min fråga om de stora transportnäten för energi .
skulle ni kunna ge ett svar på detta ?
ni oroar er över att få veta om vi skall finansiera en anläggning av kärnkraftverk någonstans med strukturfonder ? jag förenklar .
man kan säga att det inte är fråga om det .
jag har sagt er att projektvalet är medlemsstaternas sak utifrån förordningen om strukturfonderna .
kommissionens enheter är följaktligen inte systematiskt informerade om samtliga valda projekt .
ni gör dock rätt i att fråga mig , det är ert arbete och mitt är att svara .
liksom det har skett i det förflutna , måste medlemsstaterna svara då kommissionen frågar dem eller begär klargöranden .
jag skall således gå litet längre än det förtroende som vanligen delas mellan medlemsstaterna och kommissionen , och om den speciella punkt som ni nämner skall jag se efter exakt vad det handlar om .
den medlemsstat eller de berörda medlemsstaterna måste då svara mig och jag kommer genast att hänvisa svaret till er .
jag trodde mig ha svarat på frågan om de stora näten .
energisituationen varierar kraftigt beroende på område i europeiska unionen och stödet från fonderna skulle i vissa fall och för vissa områden kunna berättigas i synnerhet i de fall där anslutningen till de grundläggande energinäten ännu är underutvecklad .
det är det svar jag kan ge om bandet mellan de stora näten och strukturfonderna .
fråga nr 46 från ( h-0052 / 00 ) :
angående : strukturfonderna och additionalitetsprincipen mot bakgrund av kommissionens svar nyligen på min skriftliga fråga om strukturfonderna och additionalitetsprincipen undrar jag om kommissionen planerar att försöka ändra på reglerna om additionalitet .
skulle kommissionen ställa sig positiv till ändringar i bestämmelserna för att se till att additionalitetsprincipen gäller inte bara på medlemsstatsnivå utan även inom medlemsstater , när det gäller budgetmässiga bestämmelser för centrala regeringar och regioner eller länder som är autonoma inom en stat ?
jag skulle vilja svara maccormick att kommissionen inte planerar att ändra bestämmelserna för additionalitet , som för perioden 2000-2006 anges i artikel 11 i den allmänna förordningen för fonderna .
liksom i det förflutna anges det i dessa bestämmelser att additionalitetsprincipen skall tillämpas i förbindelsen mellan strukturfonderna och samtliga utgifter , jag säger utgifter , av medlemsstaten för utveckling .
i det avseendet måste man understryka att det är de utgifter som finansierats genom strukturfonderna som bör vara additionella .
det krävs inte att samfinansieringen av medlemsstaten skall vara det , det vill säga läggs till de befintliga utgifterna .
så länge som medlemsstaten inte minskar sina egna totala utgifter kan man anse och vi anser att strukturfonderna läggs till de nationella utgifterna och att additionalitetsprincipen således respekteras .
vad beträffar de tillämpliga budgetbestämmelserna i medlemsstaterna mellan centralregeringen och regionerna eller i de länder som har en intern självständighet , bestäms de enbart utifrån nationella överväganden och berörs således inte av additionaliteten , i enlighet med förordningarna .
jag ber om ursäkt för att ha gett detta ytterst juridiska svar .
efter kontroll är det i varje fall på det sättet som vi rättsligt och exakt i förhållande till förordningen om strukturfonderna från berlin bör definiera och förstå additionalitetsprincipen .
jag är tacksam för ett tydligt svar men naturligtvis litet besviken på dess innehåll .
vi har bara kvar artikel 11.1 som säger att anslag från fonderna får inte ersätta medlemsstaternas offentliga eller andra likvärdiga strukturella utgifter .
nåväl : det skall vara den rådande regeln .
tillåter artikel 11.1 möjligen följande praxis .
när en självstyrande region eller ett lands anslag från europeiska strukturfonderna ökar gör staten en åtföljande minskning av huvudfinansieringen till den regionen , så att det tillgängliga totala finansieringspaketet överensstämmer med en formel fastställd nationellt utan hänsyn till de strukturfondsmedel som beviljats av unionen .
är det verkligen tillåtet ?
tyvärr har jag inte tillräckligt med tid för att fördjupa mig och om herr maccormick tillåter skulle jag vilja säga honom genom att ge honom delvis rätt i hans resonemang att jag kommer att komplettera mitt svar skriftligt och åter ge honom de rättsliga grunderna både för artikel 11 i allmänhet och artikel 11.1 i synnerhet .
jag känner till , herr ledamot , med vilken kompetens ni följer alla dessa frågor .
jag känner också till de särskilda problem som finns i ert valdistrikt i skottland där vissa tvister eller diskussioner uppstår om dessa ämnen .
jag påminner dock om att på ett allmänt plan är det utgifterna från strukturfonderna som skall vara additionella , enligt alla antaganden , och det är så att så länge som medlemsstaten inte minskar sina totala utgifter läggs strukturfonderna till de nationella utgifterna och vi anser att additionalitetsprincipen respekteras .
jag skall ändå gå litet längre i mitt skriftliga svar som jag lovade er för att säga det mer objektivt och exakt .
additionalitet är också en stor fråga i wales , som jag företräder .
senast förra veckan var den en av de frågor som förde fram till ett misstroendevotum mot och avgång av förstesekreteraren i nationalförsamlingen i wales .
så sent som 1991 och 1992 vann kommissionen en strid mot förenade kungariket om additionalitet , vid tillfället kopplat till finansieringen från rechar-programmet .
detta ledde till att en överenskommelse undertecknades varmed förenade kungarikets regering lovade att införa förfaranden för att se till att eu : s medel användes för de områden som de var avsedda och var i själva verket additionella medel .
och ändå har vi fortfarande dessa problem i wales och skottland .
kan kommissionen granska denna speciella situation mot bakgrund av den överenskommelse som undertecknades med förenade kungarikets regering ?
jag förstår således , fru ledamot , att den debatt som jag hade kännedom om i skottland också pågår i wales .
jag skall kontrollera den punkt som ni anger och , om ni går med på det , kommer jag på samma gång att ge skriftligt svar på er fråga såsom jag lovade maccormick .
jag skall anstränga mig , herr talman , att ge ett kort svar genom att säga till ledamoten att den regionala utvecklingsplan som lades fram av de spanska myndigheterna den 29 oktober gör det inte möjligt för mig att dra någon slutsats om en fördelning av gemenskapens medel mellan de spanska mål 1-områdena - eftersom det handlar om i andalusien - och således de medel som var avsedda för den region som ni företräder .
jag vill således säga er , fru ledamot , att eftersom jag inte lyckades se saken klart vände jag mig till ekonomi- och finansministern , rato , med en skrivelse som jag har här från den 14 december för att be honom om vidare information om det framlagda dokumentet .
under de kommande veckorna skall kommissionen inleda förhandlingar med de spanska myndigheterna för att utarbeta gemenskapsstödramen för den nya perioden 2000-2006 och vid dessa möten , det kan jag försäkra er , kommer kommissionen att få de nödvändiga klarläggandena om fördelningen per region .
vad gäller andalusien , kommer jag således att skynda mig att meddela er personligen , om ni vill det , så snart som jag förfogar över informationen per sektor och per region .
herr kommissionär , problemet är att när aznar vänder sig till europeiska unionen för att ta betalt för samtliga andalusier , talar man om det för alla , men när aznar skall betala i form av tjänster till den regionala regeringen i andalusien , för samtliga andalusier , bortser han från fyrahundra tusen , och det är mycket allvarligt , för fyrahundra tusen barn är som om hela strasbourg , eller en större stad som granada , vore full av barn som aznar inte ser .
det är en viktig fråga och jag skulle vilja veta om herr kommissionär , för här kan man tala om barnbedrägeri , kommer att se till att andalusierna och andalusien inte luras på dessa pengar , att de pengar som europeiska unionen skall betala till andalusien mot bakgrund av folkräkningen , inbegriper de fyrahundra tusen barn som aznar inte räknar med när det gäller att förse dem med skolor och annan service .
fru ledamot , jag vill be er alla - ta inte det här som en varning - att vi bara behandlar frågor som har med gemenskapen att göra .
jag vet att dessa frågor är av stor betydelse i spanien och det finns olika visioner ...
jag kan påpeka för herr kommissionären att aznar är spaniens premiärminister .
ni kan nu besvara frågan .
fru ledamot , då jag hörde att ni har god röstkapacitet , hoppas jag att er röst var tillräckligt stark för att höras i madrid , men jag förstod att det ni sade inte var riktat direkt till mig .
jag har gett er mitt svar .
jag är angelägen om att strukturfonderna , och särskilt de som rör mål 1 , skall delas ut där det finns behov .
vi har kriterier som tillämpas och vi vet här indikativt vad varje område i europa borde eller skulle kunna få .
emellertid - jag gömmer mig inte bakom den , men jag är alltid tvungen att hänvisa till den allmänna förordningen , som jag bör diskutera med de nationella myndigheterna i varje land och med regeringen i varje land .
de har ansvaret att göra fördelningen så objektivt och rättvist som det är möjligt .
jag behöver veta i alla fall och därför sade jag att jag inte kan svara i dag .
eftersom jag inte har svaret , skrev jag till ekonomi- och finansministern den 14 december .
nu kommer den tid då jag blir otålig över att inte ha fått svar , men jag kommer att vidarebefordra det till er när jag får det .
jag beklagar att herr kommissionären än en gång har blivit delaktig i en fantasirik och i det här fallet lidelsefull inblandning .
i spanien - det vill jag påminna er alla om - befinner vi oss inte bara i valtider , det är tjugofem dagar kvar till valet .
det är en tröst för kommissionären att valen kommer att äga rum om tjugofem dagar , för sedan är det troligtvis ingen som kommer att ställa den här typen av frågor till honom längre .
jag tycker verkligen att det är viktigt att tala om att andalusien kommer att få 50 procent mer inom gemenskapens ramar och att spanien dessutom slår rekord vad gäller att förverkliga strukturfonderna , något som innebär att fördelningen sker helt i enlighet med tillämpningsbestämmelserna , att den är decentraliserad och att den ske enligt planerna för regional utveckling och de olika ramarna för gemenskapsstöd .
som en avslutning vill jag ställa en konkret fråga till herr kommissionären : anser ni att tillämpningsbestämmelserna för strukturfonderna bör ändras eller anser ni att de nuvarande fördelningskriterierna är godtagbara ?
jag tycker att debatten är mycket spännande .
jag förstår väl att den har en dimension som inte endast gäller gemenskapen .
därmed sagt att vi måste tänka på att det ständigt är val i samtliga unionens länder .
det som är mig ett nöje det är att strukturfonderna i grunden är ett diskussionsämne i grekland och i spanien .
nyss talade vi här om medborgardebatt och offentliga debatter . desto mer man talar om europa och det som europa gör för det dagliga livet , även om man grälar litet , ju bättre är det , förutsatt att man talar om det objektivt .
jag skall inte säga vad jag känner , herr ledamot , om en eventuell förändring av förordningen om strukturfonderna .
den antogs just i berlin i förra året . jag genomför den för de kommande sex åren .
vi kommer att tala om den med anledning av betänkandet om sammanhållning som är ett viktigt möte för mig här , med er , och inför er , för att göra en sammanfattning och på samma gång dra upp riktlinjer , och det ögonblick kommer i början av nästa år , då vi skall ta upp eventuella justeringar och eventuella ändringar .
jag ber er , låt mig just nu tillämpa den förordning som ännu inte tillämpats , eftersom den är daterad i berlin .
tack så mycket , herr barnier , för era svar .
frågorna 48 till 50 kommer att besvaras skriftligen .
fråga nr 51 från ( h-0049 / 00 ) :
angående : nya lokaler för byrån för harmonisering inom den inre marknaden för närvarande fortsätter byrån för harmonisering inom den inre marknaden att arbeta i sina gamla provisoriska lokaler trots att den nya byggnaden invigdes i juni 1999 . dessa ovanliga omständigheter motiverar följande fråga till kommissionen :
vilka är orsakerna till att byrån för harmonisering inom den inre marknaden ännu inte flyttat in i de nya lokalerna ?
ledamoten ställde en fråga i det här ämnet i november 1999 och jag skulle gärna vilja hänvisa till det svaret .
dessutom har jag med anledning av den nya frågan bett ordföranden för byrån för harmonisering inom den inre marknaden , alicante-byrån alltså , om en kommentar och jag kan därför för byråns räkning meddela ledamoten följande :
byrån är ännu inte klar att flytta in i den nya byggnaden .
tyvärr har vissa tidsfrister överskridits .
ett antal tekniska arbeten återstår , till exempel ett datornät , arkivutrymmen , en restaurang och möbler .
harmoniseringsbyrån håller på med detta och räknar med att flyttningen till den nya byggnaden skall kunna ske i juni .
föregående fråga föranledde oss att tala om valen .
jag tror att saken kom upp i samband med den frågan för ni , herr kommissionär , var inte med på den så illusoriskt kallade &quot; officiella invigningen &quot; av sätet för byrån för harmonisering inom den inre marknaden den 9 juni , mitt under valkampanjen , och sådana äger inte bara rum i spanien inför europavalen utan även inför de lokala och regionala valen .
om ni hade varit där , skulle ni garanterat ha tyckt att det var pinsamt .
kommissionens ordförande och några kanslichefer var visserligen på plats .
mitt under pågående valkampanj höll flera auktoriteter , alla från regeringspartiet , några anföranden som var uppenbart valfläsk och som dessutom direktsändes i tv .
synnerligen märkligt var anförandet av valencias regionalpresident som ägnade sig åt att lovorda den spanska regeringens liksom den egna regionala regeringens insatser , något som inte alls hörde till saken .
att mitt under pågående valkampanj inviga en byggnad som inte är färdig , och som åtta månader efter invigningen inte har kunnat användas , har skapat en ytterst pinsam situation för den spanska regeringen .
det bekymrar mig inte att den spanska regeringen har gjort bort sig , för när allt kommer omkring är det deras ansvar , däremot bekymrar det mig att kommissionen gör det genom att med sin närvaro garantera ett sådant icke representativt agerande .
därför vill jag fråga er , herr kommissionär : finner ni det normalt att inviga en byggnad mitt under en valkampanj innan den ens är färdig ?
finner ni det normalt att kommissionen genom sin närvaro garanterar ett sådant icke representativt agerande från den spanska regeringens sida ?
det hör inte till mina uppgifter att uttala mig om inrikespolitiska situationer i den ena eller den andra medlemsstaten .
därför vill jag heller inte kommentera den situation som berenguer nyss tog upp .
jag måste erkänna att jag inte känner till av vilken anledning en viss öppningshögtid i spanien äger rum .
jag kan dock säga att jag hoppas att den här byggnaden äntligen skall tas i bruk så snart som möjligt .
vidare vill jag tala om att jag själv hoppas att vara närvarande i alicante i slutet av maj för att tala vid en konferens där .
jag hoppas att byggnaden då skall ha tagits i bruk .
jag vill påpeka för kommissionären att det inte rör sig om en valfråga .
som medlemmar av utskottet för rättsliga frågor och den inre marknaden har vi sett hur denna institution har skapats och det är uppenbart att den invigdes av valmässiga skäl .
i dag - ett år senare - har den fortfarande inte tagits i bruk , och det innebär att kommissionen använde pengar på en falsk invigning .
man kan gott fråga sig om en användning av medel till en falsk invigning var motiverad .
ännu en gång , kommissionen håller sig inte sysselsatt med skälen till olika handlingar i medlemsstaterna .
kommissionen bryr sig om det som tillkännages offentligt och vad som görs .
vi tänker inte ge oss in i något som på franska kallas un procès d &apos; intention .
vi bryr oss om offentliga , officiella handlingar och händelser och inte eventuella bakomliggande motiv .
därför tycker jag också att det i det här fallet är svårt att svara medina på hans fråga .
kommissionen undrar inte över av vilken anledning något sker tidigare eller senare , förutom att kommissionen uppskattar att en byggnad , som för den här byrån , öppnas och tas i bruk så snabbt som möjligt .
vidare håller sig kommissionen inte heller sysselsatt med om vissa utgifter skedde reellt eller virtuellt .
för min del är alla utgifter reella .
vidare låter jag historien vara som den är .
eftersom frågeställaren är frånvarande , bortfaller fråga nr 52 .
eftersom de behandlar samma ämne , kommer frågorna 53 och 54 att tas upp tillsammans .
fråga nr 53 från ( h-0057 / 00 ) :
angående : svenska undantagsregler vad gäller införsel av alkoholhaltiga drycker över gränsen sverige har i dag ett undantag till år 2004 som medger en begränsning av alkoholhaltiga drycker över gränsen .
svenska regeringen och en stor folkopinion har uttryckt att detta undantag måste förlängas av folkhälsoskäl .
kan kommissionen redogöra för sin inställning till det svenska undantaget beträffande införsel av alkoholhaltiga drycker ?
fråga nr 54 från ( h-0117 / 00 ) :
angående : alkoholmonopol och den inre marknaden vilka åtgärder avser kommissionen att vidta för att förhindra den förlängning av det statliga alkoholmonopolet som sverige uppenbarligen planerar , och de införselrestriktioner som följer därav , samt för att se till att den inre marknadens bestämmelser får genomslag ?
jag skulle vilja besvara de här två frågorna på följande sätt .
vid tillträdet till europeiska unionen fick sverige behålla de kvantitativa begränsningarna för alkoholhaltiga drycker som resenärer får föra in i landet från andra medlemsstater .
det här undantaget från principen om fri rörlighet för varor och personer slutar att gälla den 30 juni i år .
sverige vill nu ha en förlängning av den här åtgärden i ytterligare fem år eftersom det skulle vara nödvändigt för att skydda folkhälsan .
min inställning i den här frågan är tydlig .
sverige har nu haft tillräckligt god tid på sig sedan anslutningen till unionen för att anpassa sin politik till ett tillstånd utan sådana importrestriktioner .
därför ser jag inget skäl till varför jag skulle föreslå en förlängning av det här undantaget .
europeiska medborgare har rätt att för egen räkning köpa varor inklusive skatter , i vilken medlemsstat de vill och sedan ta med dessa varor till en annan medlemsstat utan att de här varorna måste genomgå kontroller och utan att nya skatter eventuellt måste betalas .
det är en grundprincip för den inre marknaden och avvikelser från den principen måste vara undantag och tidsbegränsade .
vi vill garantera att svenska medborgare nu också skall kunna åtnjuta fördelarna med den inre marknaden , precis som andra medborgare i europeiska unionen kan göra .
det betyder inte alls att jag inte delar oron i sverige angående de möjliga hälsoproblem som kan förorsakas av alkoholmissbruk .
en undersökning som nyligen gjordes av professor lindgren vid universitetet i lund visade dock att ett avskaffande av begränsningarna inte skulle leda till en högre alkoholkonsumtion i sverige .
jag har redan vid två tillfällen kunnat diskutera min hållning med bosse ringholm , sveriges finansminister .
förra veckan diskuterade jag också den här frågan med den svenska riksdagens finansutskott .
det är nu upp till den svenska regeringen att vidta lämpliga åtgärder .
tack för svaret , herr kommissionär .
jag vill bara beklaga att det står fel i min fråga till kommissionen .
det står nämligen år 2004 , men det skall naturligtvis vara den 1 juli år 2000 .
jag har till viss del förståelse för kommissionens ståndpunkt att undantag skall vara tillfälliga .
det är en regel som är normal .
ändå skulle jag vilja ställa två frågor : tänker ni ändå ta upp fortsatta diskussioner med den svenska regeringen om en förlängning av undantagen , exempelvis så länge som danmark och finland har undantag ?
min andra fråga handlar om den samlade alkoholpolitiken .
man kan ju se detta som en fråga rörande den inre marknaden , men också som en folkhälsofråga för hela eu .
vilken roll spelar alkoholpolitiken i kommissionens arbete , och vilken roll spelar folkhälsoaspekterna ?
alkoholpolitiken i hela europa handlar inte bara om den inre marknaden , utan också om folkhälsan .
hade vi totalt sett betraktat dessa aspekter , hade det kanske varit lättare att föra diskussionen med sverige .
får jag be att få tacka herr andersson för fortsättningen på hans första fråga och den frågan vill jag svara på så här .
för det första så har finland och danmark undantag från grundregeln om fri rörlighet för varor fram till år 2003 .
de länderna håller på att vidta förberedande åtgärder så att de är klara för fri tillgång till alkoholhaltiga produkter år 2003 .
när det gäller sverige så är situationen litet annorlunda .
där beslutade man 1995 om en undantagsperiod på fem år och den går ut nu .
jag har ännu inte hört några argument som skulle kunna ligga till grund för att kommissionen borde förlänga den perioden .
för det andra så förs ständiga förhandlingar med den svenska regeringen .
jag kan meddela andersson att jag måndagen den 6 mars reser till stockholm för att där samtala med minister ringholm , med svenska riksdagsledamöter och om så önskas även med statsministern eller med andra ministrar , för att prata vidare om den här frågan som - det inser jag helt och fullt - ger anledning till starka politiska känslor i sverige .
för det tredje så förstår jag naturligtvis mycket väl att hälsoaspekten av den här frågan är viktig .
jag upprepar för andra gången att professor lindgren vid universitetet i lund har sagt att , vad som än sker med avseende på importbegränsningarna , alkoholkonsumtionen i sverige kommer att ligga kvar på samma nivå .
frågan är då naturligtvis var den mängd alkohol som inte förs in av resenärer då kommer ifrån .
svaret är att den antingen smugglas in eller också tillverkas den av svenska invånare själva och som andersson vet så är det ett mycket farligt och ohälsosamt förfarande .
andersson verkar tro att hälsosituationen går framåt om vi begränsar importen av alkohol .
i det fallet skulle inte bara sverige , utan alla länder i europeiska unionen vara tvungna att utgå från principen att all försäljning av alkohol skall förbjudas .
vi hade ett sådant exempel i förenta staterna .
andersson känner säkerligen till det som då kallades för prohibition .
han vet också vilka följder det hade för maffians verksamhet i förenta staterna , där man slutligen också gjorde slut på denna prohibition .
allt det här betyder att man naturligtvis måste skydda hälsan men inte genom att förbjuda alkohol , det hjälper nämligen inte .
herr talman ! det handlar ju i verkligheten om intäkter från det svenska alkoholmonopolet , och om den svenska regeringen säger att den måste använda dem för att täcka kostnader för hälsovården , så är detta ändå ett bevis för att det innebär en snedvridning av konkurrensen , ty andra länder måste själva finansiera sina hälsovårdskostnader , utan att förfoga över något alkoholmonopol .
min fråga gäller om ni också känner till undersökningar om att en måttlig konsumtion av alkohol av hög kvalitet , alltså exempelvis frankiskt vin eller bayerskt öl , rent av är hälsofrämjande , och att det därigenom rent av skulle ske en avlastning av den svenska statsbudgeten ?
om jag förstått det rätt så har posselt börjat peka på skatteaspekterna av den här frågan .
jag tror mig också veta att den höga skatten på alkoholhaltiga drycker i sverige har sitt ursprung år 1638 och att staten sedan dess får en ansenlig del av sina skatteinkomster från försäljningen av alkoholhaltiga produkter .
som ni vet så är det nu ett statligt monopol i sverige , vilket i sig inte heller är helt i enlighet med eu-lagstiftningen .
när det gäller alkoholens hälsosamma verkan - för jag tror att posselt talade om det också - så är jag helt ense med honom : jag tror att en bra flaska vin kan vara mycket bra för hälsan och socialt sett dessutom mycket angenäm . kanske kan posselt , andersson och jag själv träffas i parlamentets bar en dag och dricka en akvavit tillsammans .
herr talman ! jag lyssnade med intresse till kommissionärens svar på kravet att tillämpa den inre marknadens bestämmelser .
jag undrar om han kan säga om han anser sitt svar vara i överensstämmelse med kommissionens underlåtenhet att dra den franska regeringen inför eg-domstolen avseende tillämpningen av frankrikes &quot; loi et vin &quot; , som effektivt hindrar den inre marknadens bestämmelser att gälla vid försäljning av alkohol och alkoholprodukter i frankrike ?
kan vi nu förvänta oss att europeiska kommissionen vidtar åtgärder mot den franska republiken hos eg-domstolen ?
jag skulle vilja kort besvara den fråga som ställdes av ärade ledamoten eftersom detta ärende nu är under övervägande hos kommissionen .
kommissionen måste fatta ett beslut om ärendet är avslutat eller om det skall hänskjuta det till eg-domstolen .
mitt svar är kanske inte tillfredsställande just nu , men jag lovar den ärade ledamoten att kommissionen skall fatta det beslutet inom några veckor .
jag ber om ledamöternas förståelse för denna lilla försening av kommissionens beslut .
herr kommissionär ! har ni något skäl med hänsyn till folkhälsa till en skillnad i skattesats för till exempel , skotsk whisky eller franskt bordeauxvin eller mina kollegors bayerska öl ?
kan ni tänka er en likvärdig grund alkoholbeskattning i europa ?
frågan om punktskatter som den ärade ledamoten hänvisar till är den berörda medlemsstatens prerogativ .
kommissionen har inga medel att genomdriva någon särskild minskning eller ökning av punktskatter på alkoholprodukter eller några andra produkter .
mot slutet av detta år kommer kommissionen att överlämna en rapport om skillnaderna i punktskatter mellan medlemsstater .
den kommer utan tvivel att leda till diskussioner både med parlamentet och rådet om det nuvarande läget i denna fråga , vilket tyder på att det finns ganska stora skillnader i punktskattesatser mellan medlemsstater .
exempelvis , och jag tror att den ärade hänvisade till detta , tillämpas inga punktskatter på vin i frankrike medan de tillämpas i förenade kungariket .
det leder till en snedvridning av den inre marknaden eftersom vin smugglas från frankrike till förenade kungariket .
frågan gäller i synnerhet förhållandet mellan punktskatter och alkoholhalten i de varor som är punktskattepliktiga .
kommissionen har inga möjligheter att påverka i denna fråga .
i sverige används punktskatter rent av för att minska alkoholkonsumtionen .
även om detta leder till en skillnad i punktskattesats mellan sverige och andra medlemsstater i unionen - och det i sig självt ökar gränssmugglingen av alkoholprodukter - är det ett lagligt instrument för att minska alkoholkonsumtionen .
det finns naturligtvis efterfråge-elasticitet , i detta fall efterfråge-elasticitet rörande pris .
jag är inte exakt säker på vad det är men det är inte noll , därför bör den ge någon effekt .
min fråga skulle ha blivit nästan exakt den som purvis ställde , men jag skulle vilja gå vidare i frågan .
förutsatt , som ni säger , att punktskatter är medlemsstaternas prerogativ , kan ändå användning av det prerogativet på ett sätt som är diskriminerande mot producenter i en del av gemenskapen till skillnad mot andra fortfarande strida mot den inre marknadens princip .
om vi till exempel tar vad purvis och jag skulle tänka på , de maltwhiskyproducerande delarna av skotska högländerna - ett verkligt ytterområde i europa med hårda ekonomiska villkor , ett helt lantbrukssamhälle liksom ett destilleringssamhälle beroende av detta - en generell praxis att beskatta alkoholen i skotsk whisky , holländsk gin eller dansk akvavit mer än alkohol i öl eller vin tycker jag verkar diskriminerande och en diskriminerande tillämpning av något som onekligen ligger inom medlemsstaternas prerogativ .
får jag försäkra maccormick och övriga ledamöter av detta parlamentet att den nuvarande situationen med punktskatter som skiljer sig mellan medlemsstater är verkligen något som inte är bra för den inre marknadens funktion .
vi måste begränsa oss till alkoholprodukter .
om man ser på olja till exempel finner man att punktskattesatserna i tyskland skiljer sig från dem i holland och följaktligen åker holländska motorister över gränsen och tankar i tyskland .
det är i själva verket en snedvridning av den inre marknaden .
om jag fick göra som jag ville skulle jag svänga en trollstav och likställa alla punktskatter i hela europa .
följden skulle bli att smuggling upphörde utom i de fall produkter var väsentligt dyrare i en medlemsstat än i en annan .
men jag har inget trollspö och jag får inte göra som jag vill .
detta är ett område för enhällighet , som maccormick vet , och om inte alla medlemsstater går med på att likställa punktskatter , kommer det inte att ske .
ännu en gång , mot slutet av detta år kommer kommissionen att överlämna en rapport om det nuvarande läget rörande punktskatter och jag finns naturligtvis tillgänglig för diskussioner med parlamentet om den rapporten .
tack så mycket herr kommissionär .
i dag kommer vi att följa ert råd och dricka ett - eller kanske två - glas vin från alsace . vi vet inte vilka pålagor det vinet har , men jag förmodar att även det är belagt med höga skatter .
eftersom tiden för frågor till kommissionen är ute , kommer frågorna nr 55 till 114 att besvaras skriftligen .
jag förklarar härmed frågestunden med frågor till kommissionen avslutad .
( sammanträdet avbröts kl. 19.30 och återupptogs kl. 21.00 )
gemenskapsåtgärder på vattenpolitikens område ( fortsättning på debatten )
nästa punkt på föredragningslistan är fortsatt debatt om andrabehandlingsrekommendationen om gemenskapsåtgärder på vattenpolitikens område .
herr talman ! situationen för europas sötvatten är inte lika allvarlig som i andra del av världen , men rent allmänt är det ett bevisat faktum att efterfrågan på vatten ständigt ökar samtidigt som kvaliteten minskar .
därtill kommer de problem med förorening av vattnet som de potentiella nya medlemsstaterna i öst tampas med .
för övrigt har en behållare med cyanid just gått sönder i rumänien , något som utgör ett hot mot grundvattenakviferer som förser jugoslaviens befolkning med vatten .
jag har förstått det som att wallström , vars närvaro här i kväll jag uppskattar , kommer att besöka området .
jag tror inte att något land , någon regering och givetvis inte någon medlem av parlamentet kan låta bli att erkänna behovet av detta direktiv för att sätta stopp för den nuvarande uppdelningen av vattenpolitiken och underlätta igångsättandet av ett program med specifika åtgärder för olika vattendrag .
det har varit svårt och komplicerat att ta fram direktivet , det är många intressen som står på spel och åsikterna är delade .
jag tvivlar inte på att den här mandatperiodens föredragande , lienemann , har lagt ned stor möda och stort engagemang på att förena och återförena olika ståndpunkter , och hon har i stor utsträckning lyckats med det .
däremot är det nästan omöjligt att känna till och rättvist bedöma alla situationer och förväntningar .
jag kommer från ett land vars södra del vetter mot medelhavet och där tillgången till vatten historiskt sett har berott på växlingarna i ett ombytligt klimat och markens svåra beskaffenhet .
i medelhavsområdet har man varit tvungen att kämpa för sin utveckling genom att sträva efter att övervinna dessa svårigheter sekel efter sekel , år efter år , dag efter dag fram tills i dag .
som viktig betraktar vi därför direktivets praktiska tillämpning av den skyldighet som fastslås i artikel 164 i fördraget angående att i gemenskapslagstiftningen skall hänsyn tas till regionernas mångfald .
i tillämpningen av just denna princip protesterar den spanska delegationen i europeiska folkpartiet mot ändringsförslagen 4 - stycke 21 - , 13 och 49 - artikel 11d ) - , eftersom de utgör starka begränsningar på ett område som är medlemsstaternas , nämligen regleringen av vattenresurserna .
det skulle vara mycket svårt för gemenskapen att fastställa villkoren för reglerandet av dessa i de olika regionerna , med tanke på den interna balans som alltid står på spel och som under alla omständigheter kräver goda kunskaper om de olika områden och intressen som berörs .
likaså förkastar vi de ändringsförslag enligt vilka man vill inbegripa den totala vattenkostnaden år 2010 .
det råder ingen tvekan om att vi måste fastställa vattenpriser som främjar en effektiv användning , men som samtidigt gör att konkurrenskraften bevaras inom de produktiva sektorerna i de minst gynnade regionerna och inte hindrar en rättmätig utveckling .
slutligen vill jag nämna något angående ändringsförslagen om farliga ämnen , där det fastslås att en nollgradig eller nära nollgradig förgiftning skall uppnås .
hittills har ingen nollgradig förgiftning upptäckts i samband med mänskliga aktiviteter .
mina damer och herrar , vi kommer inte att göra målen i detta viktiga direktiv rättvisa om vi inte kan förse det med den flexibilitet och anpassbarhet som krävs för att garantera att direktivet uppfylls .
jag hoppas att parlamentet än en gång röstar utifrån verkligheten och med respekt för subsidiaritetsprincipen och söker uppnå en bra jämvikt mellan miljömålen och de ekonomiska och sociala hänsynen , de tre viktiga komponenterna för att uppnå en hållbar utveckling som vi alla så gärna vill ha .
herr talman , ärade kommissionär ! detta är ett mycket viktigt direktiv .
målsättningen är ju att förbättra vattenkvaliteten och säkerheten i vattenförsörjningen .
medborgarna måste ha rätt till rent vatten .
det är viktigt för såväl miljön som för folkhälsan .
jag talar inte alls för egen del , eftersom jag händelsevis råkar höra till de få lyckligt lottade européer som kan dricka vatten direkt från den egna sjön .
vi måste se till att vi snabbt kommer igång med att förbättra vattenkvaliteten .
vi måste genast börja arbeta på det .
det är viktigt att tidtabellen är ambitiös .
jag anser det inte vara för ambitiöst om vi utgår ifrån att vi år 2020 inte längre släpper ut föroreningar i vattnen och att vi strävar efter att till dess uppnå en nollnivå när det gäller föroreningar och giftiga ämnen .
det är ju fråga om att vi gör det som är tekniskt möjligt ; mer än så kan det ju inte vara frågan om , men vi måste vara tillräckligt ambitiösa .
jag vill göra er uppmärksamma på en sak som också har diskuterats tidigare .
jag anser att utskottet för miljö , folkhälsa och konsumentfrågor alltför snävt avgränsat frågan om transport av vatten .
detta är inte enbart spaniens problem , det är också de nordiska ländernas problem och jag hoppas verkligen att man i dessa frågor förlitar sig på nationella lösningar då dessa miljömässigt och ekonomiskt sett är bättre än de som nu framförs i direktivet .
herr talman , fru kommissionär ! grattis , lienemann , till ett utmärkt arbete !
vatten och luft omger oss överallt .
vi delar dem med alla människor på denna jord .
vatten är en förutsättning för mänskligt liv .
och vi blir alltfler som lever i detta liv .
schleicher antydde tidigare i dag att det skulle vara orealistiskt med rent vatten .
ingenting kan vara mer fel !
det är orealistiskt att successivt försämra vattenkvaliteten , att successivt försämra livsförutsättningarna .
särskilt orealistiskt är det för jordbruket , som är mest beroende av en ren natur och rena resurser .
därför vill jag vädja till parlamentets ledamöter att inse att hårda krav på en ren miljö innebär den största realismen på lång sikt .
herr talman ! både vi och jag personligen stöder leinemanns betänkande , de mål det uppställer och det direktiv vi diskuterar .
vi borde emellertid försöka se litet längre .
t.ex. i mitt land , herr talman , är det ett gigantiskt problem att man ändrar flodernas lopp och torrlägger sjöar med stöd av ihåliga argument och naturligtvis med stora risker både för grundvattnet och för ytvattnet .
även om vi kommer fram till vem som beslutar om sådana ingrepp , anser jag att vi behöver gemensamma och mycket stränga regler .
det stora problemet , fru kommissionär , är dock enligt min mening planeringen för att återställa grundvattenreserverna och flodernas naturliga lopp och att åter fylla sjöarna med vatten . detta måste ske under de tio år som vi planerar för .
jag anser att man måste kunna välja och finansiera sådana projekt , eftersom de kan ha en utomordentligt stor betydelse för utvecklingspolitiken .
herr talman ! här har vi något som i grunden är ett bra åtgärd .
den lägger fast uppnåbara normer grundade på subsidiaritetsprinciper och förvaltning av vattenresurser .
dess syfte med bra dricksvattenkvalitet , för djur- och växtliv , miljön och för ekonomiska ändamål är rätt .
att förhindra miljöförstöring och vattenförsämring måste vara rätt liksom möjlighet att förvalta vattenresurser vid torka och översvämning .
vi har tre olösta problem .
det första är ledning av vatten mellan vattenområden .
det är en fråga som berör mina kollegor från spanien , irland och förenade kungariket .
ändringsförslagen 4 , 49 och 87 kan inte godkännas eftersom de skulle begränsa möjligheten för ett land att leda vatten från där det finns till där det behövs , vare sig det gäller områden med torka eller städer .
för det andra måste vi ha realistiska mål , men målsättning i alla fall .
om man granskar ändringsförslag 7 till exempel , som kräver fullständigt avlägsnande av naturligt förekommande ämnen , kan ni inse att några av de uppställda målen är orealistiska .
vidare är några av målen satta till nästan noll - på engelska är det en ganska meningslös term .
vi måste granska dessa mycket noga .
konceptet att fortsätta minskningen , såsom i ändringsförslag 58 , är mycket bättre .
för det tredje tar jag upp problemet för skotsk whisky .
skotsk whisky - särskilt maltwhisky , som är den bästa - kräver vattenextraktion som används till en viss mängd och sedan återförs till vattensystemen .
en del av det slutar i flaskan och dricks upp .
vi måste se till att man i ändringsförslag 49 och 87 tar bort undantaget om att den skall utgå så att whisky kan fortsätta att drickas som &quot; high quality &quot; , vilket innebär att man för den måste använda bra , skotskt torvvatten .
det är min tredje begäran - att vi granskar noggrant dessa åtgärder innan man godkänner hela denna åtgärd .
herr talman ! först vill jag påtala det bottenlösa hyckleriet hos dem som , samtidigt som de skryter om sitt engagemang för miljön och för vattnet , gör sig skyldiga till så brottsliga handlingar som attackerna mot jugoslavien , attacker som inte bara resulterat i tusentals döda och sårade utan också lett till ekologiska katastrofer när det gäller vattenreserverna , genom att vattnet inte bara blivit obrukbart utan också utomordentligt skadligt .
i anslutning till betänkandet skulle jag också vilja säga att principen om kostnadstäckning för vattenmyndigheterna absolut inte får tillämpas så att den leder till ökad beskattning av de ekonomiskt svagaste befolkningsgrupperna eller till att de små och medelstora jordbruken slås ut på grund av de enorma kostnaderna för bevattning .
jag vill också påpeka att speciellt i områden med akut vattenbrist som i mitt land , i synnerhet på öarna , är det absolut nödvändigt att ge bidrag till investeringar i infrastruktur .
syftet är att man skall spara på vatten , inte genom prisökning utan genom att öka tillgången på vatten framför allt genom att ta till vara det regnvatten som i dag rinner bort till ingen nytta och på sin väg till havet eroderar marken med alla de problem som detta innebär .
därför stöder jag ändringsförslag 107 av vår kollega marset campos .
dessutom är det nödvändigt att ta till vara flodvattnet bättre för att garantera fortsatt liv i områden som ständigt lider brist på vatten .
slutligen vill jag säga att det är omoraliskt av rådet att , i likhet med kommissionen , påstå att det inte behövs många konkreta hänvisningar och förtydliganden , eftersom de täcks av exemplen i direktivet eller behandlas i andra delar av direktivet .
syftet är att man vill behålla ett till hälften insynsskyddat område , vilket innebär att man under den första perioden , då direktivet tillämpas slutgiltigt , kan fatta en hel del avgörande beslut till gagn för storkapitalet .
herr talman ! jag vill först och främst säga att just skyddet av vattenmiljön , både vad gäller yt- och grundvattnet , förmodligen är ett av våra allra viktigaste åtaganden .
det är det för att vi kan säkerställa tillräckliga vattenresurser , men också i hög grad för att skydda vattenresurserna mot föroreningar , så att vi även i framtiden skall få rent dricksvatten .
att ha tillgång till rent dricksvatten är en rättighet för oss alla .
jag vill gärna uttrycka ett stort erkännande av lienemanns arbete i denna fråga .
hon har utfört ett kolossalt arbete och jag vill gärna ge mitt stöd till alla lienemanns ändringsförslag , som alla förbättrar den gemensamma ståndpunkten .
och jag skall bara betona det viktigaste .
först och främst tycker jag det är viktigt att vi fastställer vissa tydliga målsättningar för vattnets tillstånd redan före en period på tio år .
jag tycker också att det är viktigt att vi utövar påtryckningar på medlemsstaterna så att de utarbetar de nödvändiga åtgärdsprogrammen snabbare än vad som uttrycks i den gemensamma ståndpunkten .
slutligen vill jag säga att jag tycker att de åtstramningar som sker med hänsyn till betalningssystemen och prisfastställandet är korrekta , så att vi som konsumenter snabbare får en effektiv användning av vattenresurserna och samtidigt ett system som kan främja uppfyllandet av de miljömål som jag tror det råder stor enighet om .
även här tycker jag att tidsfristen fram till år 2010 är en lämplig tidsfrist .
slutligen vill jag säga att jag tycker det är mycket viktigt att vi kan inleda den gradvisa reduceringen av utsläpp av farliga ämnen . att vi kan göra det gradvist , men att vi samtidigt fastställer ett slutligt mål , dvs. år 2020 , när vi förhoppningsvis är nere på obefintliga utsläppsnivåer .
om det inte är möjligt att fastställa detta som mål , är jag naturligtvis beredd att stödja det förslag som avser att vi skall nå mycket nära noll under år 2020 .
jag tycker att lienemanns förslag utgör en bra grund för vidare förhandlingar med rådet .
herr talman ! jag vill tacka föredraganden av betänkandet för ett förtjänstfullt arbete i beredningen av ett viktigt direktiv .
den andra behandlingen av vattendirektivet kommer vid en läglig tidpunkt : de skakande nyheterna från miljökatastrofen i rumänien måste utnyttjas både i dagens debatt och då man mera allmänt dryftar miljödimensionen i samband med utvidgningen av unionen .
allra först måste man hitta de skyldiga till dådet och ställa dem till svars .
cyaniden och tungmetallerna som hamnat i floden är fruktansvärda exempel på hur en vårdslös inställning till miljön kan fördärva vattendragen i tiotals år framöver .
händelsen visar att miljönormerna och inställningen till miljön i några av de länder som ansökt om eu-medlemskap ännu befinner sig ljusår från eu-nivån .
det vore också bra om unionen än en gång övervägde hur stöden till miljöprojekt skulle kunna styras för att stödja en hållbar vattenpolitik .
med tanke på förslaget till direktiv är det bekymmersamt att man under granskningarna i utskottet för miljö , folkhälsa och konsumentfrågor inte tillräckligt beaktar de oförorenade ytvattnens betydelse för de naturliga grundvattenförekomsternas utbredning .
i finland är ytvattnen mycket rena .
tillverkningen av så kallat konstgjort grundvatten är ett ekologiskt sätt att filtrera rent ytvatten som påfyllning till grundvattenreserverna .
processen kräver inga kemiska reningsverk .
direktivet får inte äventyra denna verksamhet .